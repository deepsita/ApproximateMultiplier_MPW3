magic
tech sky130A
magscale 1 2
timestamp 1635497614
<< checkpaint >>
rect -12658 -11586 596582 715522
<< locali >>
rect 239229 456943 239263 457385
rect 274005 457215 274039 457385
rect 275569 457147 275603 457385
rect 283481 456875 283515 457385
rect 377597 456807 377631 457317
rect 380909 457079 380943 457317
rect 407589 457011 407623 457317
rect 288357 336447 288391 336685
rect 277777 336311 277811 336413
rect 283205 335971 283239 336277
rect 294521 335699 294555 336413
rect 353401 336175 353435 336413
rect 378609 336175 378643 336345
rect 378701 335903 378735 336413
rect 380909 336311 380943 336413
rect 372537 335631 372571 335869
rect 378793 335835 378827 336277
rect 382289 336175 382323 336481
rect 393237 335427 393271 336005
rect 393179 335393 393271 335427
rect 402805 335359 402839 336005
rect 413109 335359 413143 335665
rect 414581 335427 414615 335597
rect 251281 333047 251315 333285
rect 302525 323595 302559 326417
rect 258123 8109 258457 8143
rect 258089 7871 258123 7973
rect 84301 4097 84577 4131
rect 84301 4063 84335 4097
rect 320741 3723 320775 3893
rect 326295 3825 326445 3859
rect 53941 3383 53975 3621
rect 320281 3519 320315 3689
rect 329941 3383 329975 3485
rect 354229 3451 354263 3689
rect 102149 3111 102183 3281
rect 354137 3179 354171 3417
rect 359565 3179 359599 3281
rect 111165 2907 111199 3077
rect 363797 2975 363831 3825
rect 535009 3383 535043 4097
<< viali >>
rect 239229 457385 239263 457419
rect 274005 457385 274039 457419
rect 274005 457181 274039 457215
rect 275569 457385 275603 457419
rect 275569 457113 275603 457147
rect 283481 457385 283515 457419
rect 239229 456909 239263 456943
rect 283481 456841 283515 456875
rect 377597 457317 377631 457351
rect 380909 457317 380943 457351
rect 380909 457045 380943 457079
rect 407589 457317 407623 457351
rect 407589 456977 407623 457011
rect 377597 456773 377631 456807
rect 288357 336685 288391 336719
rect 382289 336481 382323 336515
rect 277777 336413 277811 336447
rect 288357 336413 288391 336447
rect 294521 336413 294555 336447
rect 277777 336277 277811 336311
rect 283205 336277 283239 336311
rect 283205 335937 283239 335971
rect 353401 336413 353435 336447
rect 378701 336413 378735 336447
rect 353401 336141 353435 336175
rect 378609 336345 378643 336379
rect 378609 336141 378643 336175
rect 380909 336413 380943 336447
rect 294521 335665 294555 335699
rect 372537 335869 372571 335903
rect 378701 335869 378735 335903
rect 378793 336277 378827 336311
rect 380909 336277 380943 336311
rect 382289 336141 382323 336175
rect 378793 335801 378827 335835
rect 393237 336005 393271 336039
rect 372537 335597 372571 335631
rect 393145 335393 393179 335427
rect 402805 336005 402839 336039
rect 402805 335325 402839 335359
rect 413109 335665 413143 335699
rect 414581 335597 414615 335631
rect 414581 335393 414615 335427
rect 413109 335325 413143 335359
rect 251281 333285 251315 333319
rect 251281 333013 251315 333047
rect 302525 326417 302559 326451
rect 302525 323561 302559 323595
rect 258089 8109 258123 8143
rect 258457 8109 258491 8143
rect 258089 7973 258123 8007
rect 258089 7837 258123 7871
rect 84577 4097 84611 4131
rect 535009 4097 535043 4131
rect 84301 4029 84335 4063
rect 320741 3893 320775 3927
rect 326261 3825 326295 3859
rect 326445 3825 326479 3859
rect 363797 3825 363831 3859
rect 320281 3689 320315 3723
rect 320741 3689 320775 3723
rect 354229 3689 354263 3723
rect 53941 3621 53975 3655
rect 320281 3485 320315 3519
rect 329941 3485 329975 3519
rect 53941 3349 53975 3383
rect 329941 3349 329975 3383
rect 354137 3417 354171 3451
rect 354229 3417 354263 3451
rect 102149 3281 102183 3315
rect 354137 3145 354171 3179
rect 359565 3281 359599 3315
rect 359565 3145 359599 3179
rect 102149 3077 102183 3111
rect 111165 3077 111199 3111
rect 535009 3349 535043 3383
rect 363797 2941 363831 2975
rect 111165 2873 111199 2907
<< metal1 >>
rect 317322 700952 317328 701004
rect 317380 700992 317386 701004
rect 429838 700992 429844 701004
rect 317380 700964 429844 700992
rect 317380 700952 317386 700964
rect 429838 700952 429844 700964
rect 429896 700952 429902 701004
rect 202782 700884 202788 700936
rect 202840 700924 202846 700936
rect 331306 700924 331312 700936
rect 202840 700896 331312 700924
rect 202840 700884 202846 700896
rect 331306 700884 331312 700896
rect 331364 700884 331370 700936
rect 313182 700816 313188 700868
rect 313240 700856 313246 700868
rect 462314 700856 462320 700868
rect 313240 700828 462320 700856
rect 313240 700816 313246 700828
rect 462314 700816 462320 700828
rect 462372 700816 462378 700868
rect 315942 700748 315948 700800
rect 316000 700788 316006 700800
rect 478506 700788 478512 700800
rect 316000 700760 478512 700788
rect 316000 700748 316006 700760
rect 478506 700748 478512 700760
rect 478564 700748 478570 700800
rect 311802 700680 311808 700732
rect 311860 700720 311866 700732
rect 494790 700720 494796 700732
rect 311860 700692 494796 700720
rect 311860 700680 311866 700692
rect 494790 700680 494796 700692
rect 494848 700680 494854 700732
rect 137830 700612 137836 700664
rect 137888 700652 137894 700664
rect 336734 700652 336740 700664
rect 137888 700624 336740 700652
rect 137888 700612 137894 700624
rect 336734 700612 336740 700624
rect 336792 700612 336798 700664
rect 309042 700544 309048 700596
rect 309100 700584 309106 700596
rect 527174 700584 527180 700596
rect 309100 700556 527180 700584
rect 309100 700544 309106 700556
rect 527174 700544 527180 700556
rect 527232 700544 527238 700596
rect 105446 700476 105452 700528
rect 105504 700516 105510 700528
rect 106182 700516 106188 700528
rect 105504 700488 106188 700516
rect 105504 700476 105510 700488
rect 106182 700476 106188 700488
rect 106240 700476 106246 700528
rect 310422 700476 310428 700528
rect 310480 700516 310486 700528
rect 543458 700516 543464 700528
rect 310480 700488 543464 700516
rect 310480 700476 310486 700488
rect 543458 700476 543464 700488
rect 543516 700476 543522 700528
rect 40494 700408 40500 700460
rect 40552 700448 40558 700460
rect 41322 700448 41328 700460
rect 40552 700420 41328 700448
rect 40552 700408 40558 700420
rect 41322 700408 41328 700420
rect 41380 700408 41386 700460
rect 307662 700408 307668 700460
rect 307720 700448 307726 700460
rect 559650 700448 559656 700460
rect 307720 700420 559656 700448
rect 307720 700408 307726 700420
rect 559650 700408 559656 700420
rect 559708 700408 559714 700460
rect 72970 700340 72976 700392
rect 73028 700380 73034 700392
rect 340874 700380 340880 700392
rect 73028 700352 340880 700380
rect 73028 700340 73034 700352
rect 340874 700340 340880 700352
rect 340932 700340 340938 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 345014 700312 345020 700324
rect 8168 700284 345020 700312
rect 8168 700272 8174 700284
rect 345014 700272 345020 700284
rect 345072 700272 345078 700324
rect 320082 700204 320088 700256
rect 320140 700244 320146 700256
rect 413646 700244 413652 700256
rect 320140 700216 413652 700244
rect 320140 700204 320146 700216
rect 413646 700204 413652 700216
rect 413704 700204 413710 700256
rect 318702 700136 318708 700188
rect 318760 700176 318766 700188
rect 397454 700176 397460 700188
rect 318760 700148 397460 700176
rect 318760 700136 318766 700148
rect 397454 700136 397460 700148
rect 397512 700136 397518 700188
rect 267642 700068 267648 700120
rect 267700 700108 267706 700120
rect 327074 700108 327080 700120
rect 267700 700080 327080 700108
rect 267700 700068 267706 700080
rect 327074 700068 327080 700080
rect 327132 700068 327138 700120
rect 321462 700000 321468 700052
rect 321520 700040 321526 700052
rect 364978 700040 364984 700052
rect 321520 700012 364984 700040
rect 321520 700000 321526 700012
rect 364978 700000 364984 700012
rect 365036 700000 365042 700052
rect 324222 699932 324228 699984
rect 324280 699972 324286 699984
rect 348786 699972 348792 699984
rect 324280 699944 348792 699972
rect 324280 699932 324286 699944
rect 348786 699932 348792 699944
rect 348844 699932 348850 699984
rect 322842 699864 322848 699916
rect 322900 699904 322906 699916
rect 332502 699904 332508 699916
rect 322900 699876 332508 699904
rect 322900 699864 322906 699876
rect 332502 699864 332508 699876
rect 332560 699864 332566 699916
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 170306 699660 170312 699712
rect 170364 699700 170370 699712
rect 171042 699700 171048 699712
rect 170364 699672 171048 699700
rect 170364 699660 170370 699672
rect 171042 699660 171048 699672
rect 171100 699660 171106 699712
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 235902 699700 235908 699712
rect 235224 699672 235908 699700
rect 235224 699660 235230 699672
rect 235902 699660 235908 699672
rect 235960 699660 235966 699712
rect 300118 699660 300124 699712
rect 300176 699700 300182 699712
rect 300762 699700 300768 699712
rect 300176 699672 300768 699700
rect 300176 699660 300182 699672
rect 300762 699660 300768 699672
rect 300820 699660 300826 699712
rect 304902 696940 304908 696992
rect 304960 696980 304966 696992
rect 580166 696980 580172 696992
rect 304960 696952 580172 696980
rect 304960 696940 304966 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 306282 683136 306288 683188
rect 306340 683176 306346 683188
rect 580166 683176 580172 683188
rect 306340 683148 580172 683176
rect 306340 683136 306346 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 302142 670692 302148 670744
rect 302200 670732 302206 670744
rect 580166 670732 580172 670744
rect 302200 670704 580172 670732
rect 302200 670692 302206 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3142 656888 3148 656940
rect 3200 656928 3206 656940
rect 350534 656928 350540 656940
rect 3200 656900 350540 656928
rect 3200 656888 3206 656900
rect 350534 656888 350540 656900
rect 350592 656888 350598 656940
rect 299382 643084 299388 643136
rect 299440 643124 299446 643136
rect 580166 643124 580172 643136
rect 299440 643096 580172 643124
rect 299440 643084 299446 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 300670 630640 300676 630692
rect 300728 630680 300734 630692
rect 580166 630680 580172 630692
rect 300728 630652 580172 630680
rect 300728 630640 300734 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 2958 618264 2964 618316
rect 3016 618304 3022 618316
rect 333238 618304 333244 618316
rect 3016 618276 333244 618304
rect 3016 618264 3022 618276
rect 333238 618264 333244 618276
rect 333296 618264 333302 618316
rect 298002 616836 298008 616888
rect 298060 616876 298066 616888
rect 580166 616876 580172 616888
rect 298060 616848 580172 616876
rect 298060 616836 298066 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3326 605820 3332 605872
rect 3384 605860 3390 605872
rect 354674 605860 354680 605872
rect 3384 605832 354680 605860
rect 3384 605820 3390 605832
rect 354674 605820 354680 605832
rect 354732 605820 354738 605872
rect 295242 590656 295248 590708
rect 295300 590696 295306 590708
rect 579798 590696 579804 590708
rect 295300 590668 579804 590696
rect 295300 590656 295306 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 296622 576852 296628 576904
rect 296680 576892 296686 576904
rect 580166 576892 580172 576904
rect 296680 576864 580172 576892
rect 296680 576852 296686 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3326 565836 3332 565888
rect 3384 565876 3390 565888
rect 338758 565876 338764 565888
rect 3384 565848 338764 565876
rect 3384 565836 3390 565848
rect 338758 565836 338764 565848
rect 338816 565836 338822 565888
rect 293862 563048 293868 563100
rect 293920 563088 293926 563100
rect 579798 563088 579804 563100
rect 293920 563060 579804 563088
rect 293920 563048 293926 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 360194 553432 360200 553444
rect 3384 553404 360200 553432
rect 3384 553392 3390 553404
rect 360194 553392 360200 553404
rect 360252 553392 360258 553444
rect 289722 536800 289728 536852
rect 289780 536840 289786 536852
rect 580166 536840 580172 536852
rect 289780 536812 580172 536840
rect 289780 536800 289786 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 291102 524424 291108 524476
rect 291160 524464 291166 524476
rect 580166 524464 580172 524476
rect 291160 524436 580172 524464
rect 291160 524424 291166 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3326 514768 3332 514820
rect 3384 514808 3390 514820
rect 342898 514808 342904 514820
rect 3384 514780 342904 514808
rect 3384 514768 3390 514780
rect 342898 514768 342904 514780
rect 342956 514768 342962 514820
rect 288342 510620 288348 510672
rect 288400 510660 288406 510672
rect 580166 510660 580172 510672
rect 288400 510632 580172 510660
rect 288400 510620 288406 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3234 500964 3240 501016
rect 3292 501004 3298 501016
rect 364334 501004 364340 501016
rect 3292 500976 364340 501004
rect 3292 500964 3298 500976
rect 364334 500964 364340 500976
rect 364392 500964 364398 501016
rect 285582 484372 285588 484424
rect 285640 484412 285646 484424
rect 580166 484412 580172 484424
rect 285640 484384 580172 484412
rect 285640 484372 285646 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 286962 470568 286968 470620
rect 287020 470608 287026 470620
rect 579982 470608 579988 470620
rect 287020 470580 579988 470608
rect 287020 470568 287026 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 3510 462340 3516 462392
rect 3568 462380 3574 462392
rect 348510 462380 348516 462392
rect 3568 462352 348516 462380
rect 3568 462340 3574 462352
rect 348510 462340 348516 462352
rect 348568 462340 348574 462392
rect 154482 460844 154488 460896
rect 154540 460884 154546 460896
rect 338114 460884 338120 460896
rect 154540 460856 338120 460884
rect 154540 460844 154546 460856
rect 338114 460844 338120 460856
rect 338172 460844 338178 460896
rect 338758 460844 338764 460896
rect 338816 460884 338822 460896
rect 361758 460884 361764 460896
rect 338816 460856 361764 460884
rect 338816 460844 338822 460856
rect 361758 460844 361764 460856
rect 361816 460844 361822 460896
rect 106182 460776 106188 460828
rect 106240 460816 106246 460828
rect 339678 460816 339684 460828
rect 106240 460788 339684 460816
rect 106240 460776 106246 460788
rect 339678 460776 339684 460788
rect 339736 460776 339742 460828
rect 89622 460708 89628 460760
rect 89680 460748 89686 460760
rect 342806 460748 342812 460760
rect 89680 460720 342812 460748
rect 89680 460708 89686 460720
rect 342806 460708 342812 460720
rect 342864 460708 342870 460760
rect 342898 460708 342904 460760
rect 342956 460748 342962 460760
rect 366450 460748 366456 460760
rect 342956 460720 366456 460748
rect 342956 460708 342962 460720
rect 366450 460708 366456 460720
rect 366508 460708 366514 460760
rect 41322 460640 41328 460692
rect 41380 460680 41386 460692
rect 344370 460680 344376 460692
rect 41380 460652 344376 460680
rect 41380 460640 41386 460652
rect 344370 460640 344376 460652
rect 344428 460640 344434 460692
rect 24762 460572 24768 460624
rect 24820 460612 24826 460624
rect 347774 460612 347780 460624
rect 24820 460584 347780 460612
rect 24820 460572 24826 460584
rect 347774 460572 347780 460584
rect 347832 460572 347838 460624
rect 348510 460572 348516 460624
rect 348568 460612 348574 460624
rect 371234 460612 371240 460624
rect 348568 460584 371240 460612
rect 348568 460572 348574 460584
rect 371234 460572 371240 460584
rect 371292 460572 371298 460624
rect 3418 460504 3424 460556
rect 3476 460544 3482 460556
rect 349154 460544 349160 460556
rect 3476 460516 349160 460544
rect 3476 460504 3482 460516
rect 349154 460504 349160 460516
rect 349212 460504 349218 460556
rect 3602 460436 3608 460488
rect 3660 460476 3666 460488
rect 352282 460476 352288 460488
rect 3660 460448 352288 460476
rect 3660 460436 3666 460448
rect 352282 460436 352288 460448
rect 352340 460436 352346 460488
rect 3694 460368 3700 460420
rect 3752 460408 3758 460420
rect 353846 460408 353852 460420
rect 3752 460380 353852 460408
rect 3752 460368 3758 460380
rect 353846 460368 353852 460380
rect 353904 460368 353910 460420
rect 3786 460300 3792 460352
rect 3844 460340 3850 460352
rect 358814 460340 358820 460352
rect 3844 460312 358820 460340
rect 3844 460300 3850 460312
rect 358814 460300 358820 460312
rect 358872 460300 358878 460352
rect 3878 460232 3884 460284
rect 3936 460272 3942 460284
rect 363322 460272 363328 460284
rect 3936 460244 363328 460272
rect 3936 460232 3942 460244
rect 363322 460232 363328 460244
rect 363380 460232 363386 460284
rect 3970 460164 3976 460216
rect 4028 460204 4034 460216
rect 368106 460204 368112 460216
rect 4028 460176 368112 460204
rect 4028 460164 4034 460176
rect 368106 460164 368112 460176
rect 368164 460164 368170 460216
rect 171042 460096 171048 460148
rect 171100 460136 171106 460148
rect 334894 460136 334900 460148
rect 171100 460108 334900 460136
rect 171100 460096 171106 460108
rect 334894 460096 334900 460108
rect 334952 460096 334958 460148
rect 219342 460028 219348 460080
rect 219400 460068 219406 460080
rect 219400 460040 333192 460068
rect 219400 460028 219406 460040
rect 235902 459960 235908 460012
rect 235960 460000 235966 460012
rect 330202 460000 330208 460012
rect 235960 459972 330208 460000
rect 235960 459960 235966 459972
rect 330202 459960 330208 459972
rect 330260 459960 330266 460012
rect 333164 460000 333192 460040
rect 333238 460028 333244 460080
rect 333296 460068 333302 460080
rect 356974 460068 356980 460080
rect 333296 460040 356980 460068
rect 333296 460028 333302 460040
rect 356974 460028 356980 460040
rect 357032 460028 357038 460080
rect 333330 460000 333336 460012
rect 333164 459972 333336 460000
rect 333330 459960 333336 459972
rect 333388 459960 333394 460012
rect 284202 459892 284208 459944
rect 284260 459932 284266 459944
rect 328546 459932 328552 459944
rect 284260 459904 328552 459932
rect 284260 459892 284266 459904
rect 328546 459892 328552 459904
rect 328604 459892 328610 459944
rect 325694 459864 325700 459876
rect 316006 459836 325700 459864
rect 300762 459756 300768 459808
rect 300820 459796 300826 459808
rect 316006 459796 316034 459836
rect 325694 459824 325700 459836
rect 325752 459824 325758 459876
rect 300820 459768 316034 459796
rect 300820 459756 300826 459768
rect 281442 459688 281448 459740
rect 281500 459728 281506 459740
rect 281500 459700 287054 459728
rect 281500 459688 281506 459700
rect 285030 459620 285036 459672
rect 285088 459660 285094 459672
rect 285582 459660 285588 459672
rect 285088 459632 285588 459660
rect 285088 459620 285094 459632
rect 285582 459620 285588 459632
rect 285640 459620 285646 459672
rect 287026 459660 287054 459700
rect 292942 459688 292948 459740
rect 293000 459728 293006 459740
rect 293862 459728 293868 459740
rect 293000 459700 293868 459728
rect 293000 459688 293006 459700
rect 293862 459688 293868 459700
rect 293920 459688 293926 459740
rect 294506 459688 294512 459740
rect 294564 459728 294570 459740
rect 295242 459728 295248 459740
rect 294564 459700 295248 459728
rect 294564 459688 294570 459700
rect 295242 459688 295248 459700
rect 295300 459688 295306 459740
rect 296070 459688 296076 459740
rect 296128 459728 296134 459740
rect 296622 459728 296628 459740
rect 296128 459700 296628 459728
rect 296128 459688 296134 459700
rect 296622 459688 296628 459700
rect 296680 459688 296686 459740
rect 303982 459688 303988 459740
rect 304040 459728 304046 459740
rect 304902 459728 304908 459740
rect 304040 459700 304908 459728
rect 304040 459688 304046 459700
rect 304902 459688 304908 459700
rect 304960 459688 304966 459740
rect 305546 459688 305552 459740
rect 305604 459728 305610 459740
rect 306282 459728 306288 459740
rect 305604 459700 306288 459728
rect 305604 459688 305610 459700
rect 306282 459688 306288 459700
rect 306340 459688 306346 459740
rect 307110 459688 307116 459740
rect 307168 459728 307174 459740
rect 307662 459728 307668 459740
rect 307168 459700 307668 459728
rect 307168 459688 307174 459700
rect 307662 459688 307668 459700
rect 307720 459688 307726 459740
rect 315022 459688 315028 459740
rect 315080 459728 315086 459740
rect 315942 459728 315948 459740
rect 315080 459700 315948 459728
rect 315080 459688 315086 459700
rect 315942 459688 315948 459700
rect 316000 459688 316006 459740
rect 316586 459688 316592 459740
rect 316644 459728 316650 459740
rect 317322 459728 317328 459740
rect 316644 459700 317328 459728
rect 316644 459688 316650 459700
rect 317322 459688 317328 459700
rect 317380 459688 317386 459740
rect 318150 459688 318156 459740
rect 318208 459728 318214 459740
rect 318702 459728 318708 459740
rect 318208 459700 318708 459728
rect 318208 459688 318214 459700
rect 318702 459688 318708 459700
rect 318760 459688 318766 459740
rect 556798 459660 556804 459672
rect 287026 459632 556804 459660
rect 556798 459620 556804 459632
rect 556856 459620 556862 459672
rect 272334 459552 272340 459604
rect 272392 459592 272398 459604
rect 555418 459592 555424 459604
rect 272392 459564 555424 459592
rect 272392 459552 272398 459564
rect 555418 459552 555424 459564
rect 555476 459552 555482 459604
rect 255038 458804 255044 458856
rect 255096 458844 255102 458856
rect 580258 458844 580264 458856
rect 255096 458816 580264 458844
rect 255096 458804 255102 458816
rect 580258 458804 580264 458816
rect 580316 458804 580322 458856
rect 278682 458668 278688 458720
rect 278740 458708 278746 458720
rect 418798 458708 418804 458720
rect 278740 458680 418804 458708
rect 278740 458668 278746 458680
rect 418798 458668 418804 458680
rect 418856 458668 418862 458720
rect 280062 458600 280068 458652
rect 280120 458640 280126 458652
rect 428458 458640 428464 458652
rect 280120 458612 428464 458640
rect 280120 458600 280126 458612
rect 428458 458600 428464 458612
rect 428516 458600 428522 458652
rect 228358 458532 228364 458584
rect 228416 458572 228422 458584
rect 379146 458572 379152 458584
rect 228416 458544 379152 458572
rect 228416 458532 228422 458544
rect 379146 458532 379152 458544
rect 379204 458532 379210 458584
rect 270402 458464 270408 458516
rect 270460 458504 270466 458516
rect 421650 458504 421656 458516
rect 270460 458476 421656 458504
rect 270460 458464 270466 458476
rect 421650 458464 421656 458476
rect 421708 458464 421714 458516
rect 222838 458396 222844 458448
rect 222896 458436 222902 458448
rect 375926 458436 375932 458448
rect 222896 458408 375932 458436
rect 222896 458396 222902 458408
rect 375926 458396 375932 458408
rect 375984 458396 375990 458448
rect 277026 458328 277032 458380
rect 277084 458368 277090 458380
rect 429838 458368 429844 458380
rect 277084 458340 429844 458368
rect 277084 458328 277090 458340
rect 429838 458328 429844 458340
rect 429896 458328 429902 458380
rect 232590 458260 232596 458312
rect 232648 458300 232654 458312
rect 391934 458300 391940 458312
rect 232648 458272 391940 458300
rect 232648 458260 232654 458272
rect 391934 458260 391940 458272
rect 391992 458260 391998 458312
rect 3418 458192 3424 458244
rect 3476 458232 3482 458244
rect 373120 458232 373126 458244
rect 3476 458204 373126 458232
rect 3476 458192 3482 458204
rect 373120 458192 373126 458204
rect 373178 458192 373184 458244
rect 233878 457376 233884 457428
rect 233936 457416 233942 457428
rect 239214 457416 239220 457428
rect 233936 457388 238754 457416
rect 239175 457388 239220 457416
rect 233936 457376 233942 457388
rect 238726 457348 238754 457388
rect 239214 457376 239220 457388
rect 239272 457376 239278 457428
rect 273990 457416 273996 457428
rect 273951 457388 273996 457416
rect 273990 457376 273996 457388
rect 274048 457376 274054 457428
rect 275554 457416 275560 457428
rect 275515 457388 275560 457416
rect 275554 457376 275560 457388
rect 275612 457376 275618 457428
rect 283466 457416 283472 457428
rect 283427 457388 283472 457416
rect 283466 457376 283472 457388
rect 283524 457376 283530 457428
rect 369854 457348 369860 457360
rect 238726 457320 369860 457348
rect 369854 457308 369860 457320
rect 369912 457308 369918 457360
rect 374362 457348 374368 457360
rect 373966 457320 374368 457348
rect 231118 457240 231124 457292
rect 231176 457280 231182 457292
rect 373966 457280 373994 457320
rect 374362 457308 374368 457320
rect 374420 457308 374426 457360
rect 377582 457348 377588 457360
rect 377543 457320 377588 457348
rect 377582 457308 377588 457320
rect 377640 457308 377646 457360
rect 380894 457348 380900 457360
rect 380855 457320 380900 457348
rect 380894 457308 380900 457320
rect 380952 457308 380958 457360
rect 407574 457348 407580 457360
rect 407535 457320 407580 457348
rect 407574 457308 407580 457320
rect 407632 457308 407638 457360
rect 231176 457252 373994 457280
rect 231176 457240 231182 457252
rect 273993 457215 274051 457221
rect 273993 457181 274005 457215
rect 274039 457212 274051 457215
rect 417418 457212 417424 457224
rect 274039 457184 417424 457212
rect 274039 457181 274051 457184
rect 273993 457175 274051 457181
rect 417418 457172 417424 457184
rect 417476 457172 417482 457224
rect 275557 457147 275615 457153
rect 275557 457113 275569 457147
rect 275603 457144 275615 457147
rect 425698 457144 425704 457156
rect 275603 457116 425704 457144
rect 275603 457113 275615 457116
rect 275557 457107 275615 457113
rect 425698 457104 425704 457116
rect 425756 457104 425762 457156
rect 224218 457036 224224 457088
rect 224276 457076 224282 457088
rect 380897 457079 380955 457085
rect 380897 457076 380909 457079
rect 224276 457048 380909 457076
rect 224276 457036 224282 457048
rect 380897 457045 380909 457048
rect 380943 457045 380955 457079
rect 380897 457039 380955 457045
rect 226978 456968 226984 457020
rect 227036 457008 227042 457020
rect 407577 457011 407635 457017
rect 407577 457008 407589 457011
rect 227036 456980 407589 457008
rect 227036 456968 227042 456980
rect 407577 456977 407589 456980
rect 407623 456977 407635 457011
rect 407577 456971 407635 456977
rect 239217 456943 239275 456949
rect 239217 456909 239229 456943
rect 239263 456940 239275 456943
rect 431218 456940 431224 456952
rect 239263 456912 431224 456940
rect 239263 456909 239275 456912
rect 239217 456903 239275 456909
rect 431218 456900 431224 456912
rect 431276 456900 431282 456952
rect 283469 456875 283527 456881
rect 283469 456841 283481 456875
rect 283515 456872 283527 456875
rect 579798 456872 579804 456884
rect 283515 456844 579804 456872
rect 283515 456841 283527 456844
rect 283469 456835 283527 456841
rect 579798 456832 579804 456844
rect 579856 456832 579862 456884
rect 4798 456764 4804 456816
rect 4856 456804 4862 456816
rect 377585 456807 377643 456813
rect 377585 456804 377597 456807
rect 4856 456776 377597 456804
rect 4856 456764 4862 456776
rect 377585 456773 377597 456776
rect 377631 456773 377643 456807
rect 377585 456767 377643 456773
rect 3326 449828 3332 449880
rect 3384 449868 3390 449880
rect 233878 449868 233884 449880
rect 3384 449840 233884 449868
rect 3384 449828 3390 449840
rect 233878 449828 233884 449840
rect 233936 449828 233942 449880
rect 428458 431876 428464 431928
rect 428516 431916 428522 431928
rect 580166 431916 580172 431928
rect 428516 431888 580172 431916
rect 428516 431876 428522 431888
rect 580166 431876 580172 431888
rect 580224 431876 580230 431928
rect 556798 419432 556804 419484
rect 556856 419472 556862 419484
rect 580166 419472 580172 419484
rect 556856 419444 580172 419472
rect 556856 419432 556862 419444
rect 580166 419432 580172 419444
rect 580224 419432 580230 419484
rect 3418 411204 3424 411256
rect 3476 411244 3482 411256
rect 222838 411244 222844 411256
rect 3476 411216 222844 411244
rect 3476 411204 3482 411216
rect 222838 411204 222844 411216
rect 222896 411204 222902 411256
rect 418798 405628 418804 405680
rect 418856 405668 418862 405680
rect 579614 405668 579620 405680
rect 418856 405640 579620 405668
rect 418856 405628 418862 405640
rect 579614 405628 579620 405640
rect 579672 405628 579678 405680
rect 3234 398760 3240 398812
rect 3292 398800 3298 398812
rect 231118 398800 231124 398812
rect 3292 398772 231124 398800
rect 3292 398760 3298 398772
rect 231118 398760 231124 398772
rect 231176 398760 231182 398812
rect 425698 379448 425704 379500
rect 425756 379488 425762 379500
rect 580166 379488 580172 379500
rect 425756 379460 580172 379488
rect 425756 379448 425762 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 2774 371424 2780 371476
rect 2832 371464 2838 371476
rect 4798 371464 4804 371476
rect 2832 371436 4804 371464
rect 2832 371424 2838 371436
rect 4798 371424 4804 371436
rect 4856 371424 4862 371476
rect 429838 365644 429844 365696
rect 429896 365684 429902 365696
rect 580166 365684 580172 365696
rect 429896 365656 580172 365684
rect 429896 365644 429902 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 3326 358708 3332 358760
rect 3384 358748 3390 358760
rect 224218 358748 224224 358760
rect 3384 358720 224224 358748
rect 3384 358708 3390 358720
rect 224218 358708 224224 358720
rect 224276 358708 224282 358760
rect 417418 353200 417424 353252
rect 417476 353240 417482 353252
rect 580166 353240 580172 353252
rect 417476 353212 580172 353240
rect 417476 353200 417482 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 3142 346332 3148 346384
rect 3200 346372 3206 346384
rect 228358 346372 228364 346384
rect 3200 346344 228364 346372
rect 3200 346332 3206 346344
rect 228358 346332 228364 346344
rect 228416 346332 228422 346384
rect 220078 336676 220084 336728
rect 220136 336716 220142 336728
rect 288345 336719 288403 336725
rect 288345 336716 288357 336719
rect 220136 336688 288357 336716
rect 220136 336676 220142 336688
rect 288345 336685 288357 336688
rect 288391 336685 288403 336719
rect 288345 336679 288403 336685
rect 288434 336676 288440 336728
rect 288492 336716 288498 336728
rect 289814 336716 289820 336728
rect 288492 336688 289820 336716
rect 288492 336676 288498 336688
rect 289814 336676 289820 336688
rect 289872 336676 289878 336728
rect 291562 336676 291568 336728
rect 291620 336716 291626 336728
rect 292942 336716 292948 336728
rect 291620 336688 292948 336716
rect 291620 336676 291626 336688
rect 292942 336676 292948 336688
rect 293000 336676 293006 336728
rect 300486 336676 300492 336728
rect 300544 336716 300550 336728
rect 301314 336716 301320 336728
rect 300544 336688 301320 336716
rect 300544 336676 300550 336688
rect 301314 336676 301320 336688
rect 301372 336676 301378 336728
rect 304902 336676 304908 336728
rect 304960 336716 304966 336728
rect 328546 336716 328552 336728
rect 304960 336688 328552 336716
rect 304960 336676 304966 336688
rect 328546 336676 328552 336688
rect 328604 336676 328610 336728
rect 339494 336676 339500 336728
rect 339552 336716 339558 336728
rect 339770 336716 339776 336728
rect 339552 336688 339776 336716
rect 339552 336676 339558 336688
rect 339770 336676 339776 336688
rect 339828 336676 339834 336728
rect 342714 336676 342720 336728
rect 342772 336716 342778 336728
rect 343450 336716 343456 336728
rect 342772 336688 343456 336716
rect 342772 336676 342778 336688
rect 343450 336676 343456 336688
rect 343508 336676 343514 336728
rect 343542 336676 343548 336728
rect 343600 336716 343606 336728
rect 344278 336716 344284 336728
rect 343600 336688 344284 336716
rect 343600 336676 343606 336688
rect 344278 336676 344284 336688
rect 344336 336676 344342 336728
rect 347038 336676 347044 336728
rect 347096 336716 347102 336728
rect 347590 336716 347596 336728
rect 347096 336688 347596 336716
rect 347096 336676 347102 336688
rect 347590 336676 347596 336688
rect 347648 336676 347654 336728
rect 354030 336676 354036 336728
rect 354088 336716 354094 336728
rect 354490 336716 354496 336728
rect 354088 336688 354496 336716
rect 354088 336676 354094 336688
rect 354490 336676 354496 336688
rect 354548 336676 354554 336728
rect 355042 336676 355048 336728
rect 355100 336716 355106 336728
rect 355778 336716 355784 336728
rect 355100 336688 355784 336716
rect 355100 336676 355106 336688
rect 355778 336676 355784 336688
rect 355836 336676 355842 336728
rect 356514 336676 356520 336728
rect 356572 336716 356578 336728
rect 357158 336716 357164 336728
rect 356572 336688 357164 336716
rect 356572 336676 356578 336688
rect 357158 336676 357164 336688
rect 357216 336676 357222 336728
rect 357986 336676 357992 336728
rect 358044 336716 358050 336728
rect 358722 336716 358728 336728
rect 358044 336688 358728 336716
rect 358044 336676 358050 336688
rect 358722 336676 358728 336688
rect 358780 336676 358786 336728
rect 359458 336676 359464 336728
rect 359516 336716 359522 336728
rect 359918 336716 359924 336728
rect 359516 336688 359924 336716
rect 359516 336676 359522 336688
rect 359918 336676 359924 336688
rect 359976 336676 359982 336728
rect 360930 336676 360936 336728
rect 360988 336716 360994 336728
rect 361390 336716 361396 336728
rect 360988 336688 361396 336716
rect 360988 336676 360994 336688
rect 361390 336676 361396 336688
rect 361448 336676 361454 336728
rect 362586 336676 362592 336728
rect 362644 336716 362650 336728
rect 362862 336716 362868 336728
rect 362644 336688 362868 336716
rect 362644 336676 362650 336688
rect 362862 336676 362868 336688
rect 362920 336676 362926 336728
rect 363506 336676 363512 336728
rect 363564 336716 363570 336728
rect 364242 336716 364248 336728
rect 363564 336688 364248 336716
rect 363564 336676 363570 336688
rect 364242 336676 364248 336688
rect 364300 336676 364306 336728
rect 370406 336676 370412 336728
rect 370464 336716 370470 336728
rect 435358 336716 435364 336728
rect 370464 336688 435364 336716
rect 370464 336676 370470 336688
rect 435358 336676 435364 336688
rect 435416 336676 435422 336728
rect 215938 336608 215944 336660
rect 215996 336648 216002 336660
rect 292206 336648 292212 336660
rect 215996 336620 292212 336648
rect 215996 336608 216002 336620
rect 292206 336608 292212 336620
rect 292264 336608 292270 336660
rect 292482 336608 292488 336660
rect 292540 336648 292546 336660
rect 295426 336648 295432 336660
rect 292540 336620 295432 336648
rect 292540 336608 292546 336620
rect 295426 336608 295432 336620
rect 295484 336608 295490 336660
rect 296530 336608 296536 336660
rect 296588 336648 296594 336660
rect 296898 336648 296904 336660
rect 296588 336620 296904 336648
rect 296588 336608 296594 336620
rect 296898 336608 296904 336620
rect 296956 336608 296962 336660
rect 300762 336608 300768 336660
rect 300820 336648 300826 336660
rect 327534 336648 327540 336660
rect 300820 336620 327540 336648
rect 300820 336608 300826 336620
rect 327534 336608 327540 336620
rect 327592 336608 327598 336660
rect 341242 336608 341248 336660
rect 341300 336648 341306 336660
rect 342438 336648 342444 336660
rect 341300 336620 342444 336648
rect 341300 336608 341306 336620
rect 342438 336608 342444 336620
rect 342496 336608 342502 336660
rect 349614 336608 349620 336660
rect 349672 336648 349678 336660
rect 353938 336648 353944 336660
rect 349672 336620 353944 336648
rect 349672 336608 349678 336620
rect 353938 336608 353944 336620
rect 353996 336608 354002 336660
rect 355686 336608 355692 336660
rect 355744 336648 355750 336660
rect 355962 336648 355968 336660
rect 355744 336620 355968 336648
rect 355744 336608 355750 336620
rect 355962 336608 355968 336620
rect 356020 336608 356026 336660
rect 359090 336608 359096 336660
rect 359148 336648 359154 336660
rect 360010 336648 360016 336660
rect 359148 336620 360016 336648
rect 359148 336608 359154 336620
rect 360010 336608 360016 336620
rect 360068 336608 360074 336660
rect 362034 336608 362040 336660
rect 362092 336648 362098 336660
rect 362678 336648 362684 336660
rect 362092 336620 362684 336648
rect 362092 336608 362098 336620
rect 362678 336608 362684 336620
rect 362736 336608 362742 336660
rect 369762 336608 369768 336660
rect 369820 336648 369826 336660
rect 436094 336648 436100 336660
rect 369820 336620 436100 336648
rect 369820 336608 369826 336620
rect 436094 336608 436100 336620
rect 436152 336608 436158 336660
rect 214558 336540 214564 336592
rect 214616 336580 214622 336592
rect 293310 336580 293316 336592
rect 214616 336552 293316 336580
rect 214616 336540 214622 336552
rect 293310 336540 293316 336552
rect 293368 336540 293374 336592
rect 296622 336540 296628 336592
rect 296680 336580 296686 336592
rect 326154 336580 326160 336592
rect 296680 336552 326160 336580
rect 296680 336540 296686 336552
rect 326154 336540 326160 336552
rect 326212 336540 326218 336592
rect 345566 336540 345572 336592
rect 345624 336580 345630 336592
rect 349798 336580 349804 336592
rect 345624 336552 349804 336580
rect 345624 336540 345630 336552
rect 349798 336540 349804 336552
rect 349856 336540 349862 336592
rect 372246 336540 372252 336592
rect 372304 336580 372310 336592
rect 442994 336580 443000 336592
rect 372304 336552 443000 336580
rect 372304 336540 372310 336552
rect 442994 336540 443000 336552
rect 443052 336540 443058 336592
rect 209038 336472 209044 336524
rect 209096 336512 209102 336524
rect 296714 336512 296720 336524
rect 209096 336484 296720 336512
rect 209096 336472 209102 336484
rect 296714 336472 296720 336484
rect 296772 336472 296778 336524
rect 299382 336472 299388 336524
rect 299440 336512 299446 336524
rect 327074 336512 327080 336524
rect 299440 336484 327080 336512
rect 299440 336472 299446 336484
rect 327074 336472 327080 336484
rect 327132 336472 327138 336524
rect 329098 336472 329104 336524
rect 329156 336512 329162 336524
rect 333974 336512 333980 336524
rect 329156 336484 333980 336512
rect 329156 336472 329162 336484
rect 333974 336472 333980 336484
rect 334032 336472 334038 336524
rect 348510 336472 348516 336524
rect 348568 336512 348574 336524
rect 363598 336512 363604 336524
rect 348568 336484 363604 336512
rect 348568 336472 348574 336484
rect 363598 336472 363604 336484
rect 363656 336472 363662 336524
rect 373350 336472 373356 336524
rect 373408 336512 373414 336524
rect 373902 336512 373908 336524
rect 373408 336484 373908 336512
rect 373408 336472 373414 336484
rect 373902 336472 373908 336484
rect 373960 336472 373966 336524
rect 374822 336472 374828 336524
rect 374880 336512 374886 336524
rect 375190 336512 375196 336524
rect 374880 336484 375196 336512
rect 374880 336472 374886 336484
rect 375190 336472 375196 336484
rect 375248 336472 375254 336524
rect 375926 336472 375932 336524
rect 375984 336512 375990 336524
rect 376662 336512 376668 336524
rect 375984 336484 376668 336512
rect 375984 336472 375990 336484
rect 376662 336472 376668 336484
rect 376720 336472 376726 336524
rect 377030 336472 377036 336524
rect 377088 336512 377094 336524
rect 377858 336512 377864 336524
rect 377088 336484 377864 336512
rect 377088 336472 377094 336484
rect 377858 336472 377864 336484
rect 377916 336472 377922 336524
rect 380250 336472 380256 336524
rect 380308 336512 380314 336524
rect 380710 336512 380716 336524
rect 380308 336484 380716 336512
rect 380308 336472 380314 336484
rect 380710 336472 380716 336484
rect 380768 336472 380774 336524
rect 381998 336472 382004 336524
rect 382056 336512 382062 336524
rect 382182 336512 382188 336524
rect 382056 336484 382188 336512
rect 382056 336472 382062 336484
rect 382182 336472 382188 336484
rect 382240 336472 382246 336524
rect 382277 336515 382335 336521
rect 382277 336481 382289 336515
rect 382323 336512 382335 336515
rect 449894 336512 449900 336524
rect 382323 336484 449900 336512
rect 382323 336481 382335 336484
rect 382277 336475 382335 336481
rect 449894 336472 449900 336484
rect 449952 336472 449958 336524
rect 125502 336404 125508 336456
rect 125560 336444 125566 336456
rect 125560 336416 270586 336444
rect 125560 336404 125566 336416
rect 114462 336336 114468 336388
rect 114520 336376 114526 336388
rect 269942 336376 269948 336388
rect 114520 336348 269948 336376
rect 114520 336336 114526 336348
rect 269942 336336 269948 336348
rect 270000 336336 270006 336388
rect 270558 336376 270586 336416
rect 271782 336404 271788 336456
rect 271840 336444 271846 336456
rect 272794 336444 272800 336456
rect 271840 336416 272800 336444
rect 271840 336404 271846 336416
rect 272794 336404 272800 336416
rect 272852 336404 272858 336456
rect 276014 336404 276020 336456
rect 276072 336444 276078 336456
rect 277765 336447 277823 336453
rect 277765 336444 277777 336447
rect 276072 336416 277777 336444
rect 276072 336404 276078 336416
rect 277765 336413 277777 336416
rect 277811 336413 277823 336447
rect 277765 336407 277823 336413
rect 277854 336404 277860 336456
rect 277912 336444 277918 336456
rect 279786 336444 279792 336456
rect 277912 336416 279792 336444
rect 277912 336404 277918 336416
rect 279786 336404 279792 336416
rect 279844 336404 279850 336456
rect 282638 336404 282644 336456
rect 282696 336444 282702 336456
rect 283374 336444 283380 336456
rect 282696 336416 283380 336444
rect 282696 336404 282702 336416
rect 283374 336404 283380 336416
rect 283432 336404 283438 336456
rect 288345 336447 288403 336453
rect 288345 336413 288357 336447
rect 288391 336444 288403 336447
rect 294414 336444 294420 336456
rect 288391 336416 294420 336444
rect 288391 336413 288403 336416
rect 288345 336407 288403 336413
rect 294414 336404 294420 336416
rect 294472 336404 294478 336456
rect 294509 336447 294567 336453
rect 294509 336413 294521 336447
rect 294555 336444 294567 336447
rect 323578 336444 323584 336456
rect 294555 336416 323584 336444
rect 294555 336413 294567 336416
rect 294509 336407 294567 336413
rect 323578 336404 323584 336416
rect 323636 336404 323642 336456
rect 347406 336404 347412 336456
rect 347464 336444 347470 336456
rect 353389 336447 353447 336453
rect 353389 336444 353401 336447
rect 347464 336416 353401 336444
rect 347464 336404 347470 336416
rect 353389 336413 353401 336416
rect 353435 336413 353447 336447
rect 353389 336407 353447 336413
rect 367830 336404 367836 336456
rect 367888 336444 367894 336456
rect 378689 336447 378747 336453
rect 378689 336444 378701 336447
rect 367888 336416 378701 336444
rect 367888 336404 367894 336416
rect 378689 336413 378701 336416
rect 378735 336413 378747 336447
rect 378689 336407 378747 336413
rect 379882 336404 379888 336456
rect 379940 336444 379946 336456
rect 380618 336444 380624 336456
rect 379940 336416 380624 336444
rect 379940 336404 379946 336416
rect 380618 336404 380624 336416
rect 380676 336404 380682 336456
rect 380897 336447 380955 336453
rect 380897 336413 380909 336447
rect 380943 336444 380955 336447
rect 456794 336444 456800 336456
rect 380943 336416 456800 336444
rect 380943 336413 380955 336416
rect 380897 336407 380955 336413
rect 456794 336404 456800 336416
rect 456852 336404 456858 336456
rect 273254 336376 273260 336388
rect 270558 336348 273260 336376
rect 273254 336336 273260 336348
rect 273312 336336 273318 336388
rect 277302 336336 277308 336388
rect 277360 336376 277366 336388
rect 319898 336376 319904 336388
rect 277360 336348 319904 336376
rect 277360 336336 277366 336348
rect 319898 336336 319904 336348
rect 319956 336336 319962 336388
rect 347682 336336 347688 336388
rect 347740 336376 347746 336388
rect 348418 336376 348424 336388
rect 347740 336348 348424 336376
rect 347740 336336 347746 336348
rect 348418 336336 348424 336348
rect 348476 336336 348482 336388
rect 354398 336336 354404 336388
rect 354456 336376 354462 336388
rect 370498 336376 370504 336388
rect 354456 336348 370504 336376
rect 354456 336336 354462 336348
rect 370498 336336 370504 336348
rect 370556 336336 370562 336388
rect 374454 336336 374460 336388
rect 374512 336376 374518 336388
rect 378597 336379 378655 336385
rect 378597 336376 378609 336379
rect 374512 336348 378609 336376
rect 374512 336336 374518 336348
rect 378597 336345 378609 336348
rect 378643 336345 378655 336379
rect 378597 336339 378655 336345
rect 378870 336336 378876 336388
rect 378928 336376 378934 336388
rect 465074 336376 465080 336388
rect 378928 336348 465080 336376
rect 378928 336336 378934 336348
rect 465074 336336 465080 336348
rect 465132 336336 465138 336388
rect 107562 336268 107568 336320
rect 107620 336308 107626 336320
rect 267826 336308 267832 336320
rect 107620 336280 267832 336308
rect 107620 336268 107626 336280
rect 267826 336268 267832 336280
rect 267884 336268 267890 336320
rect 277765 336311 277823 336317
rect 277765 336277 277777 336311
rect 277811 336308 277823 336311
rect 279050 336308 279056 336320
rect 277811 336280 279056 336308
rect 277811 336277 277823 336280
rect 277765 336271 277823 336277
rect 279050 336268 279056 336280
rect 279108 336268 279114 336320
rect 282178 336268 282184 336320
rect 282236 336308 282242 336320
rect 283098 336308 283104 336320
rect 282236 336280 283104 336308
rect 282236 336268 282242 336280
rect 283098 336268 283104 336280
rect 283156 336268 283162 336320
rect 283193 336311 283251 336317
rect 283193 336277 283205 336311
rect 283239 336308 283251 336311
rect 321554 336308 321560 336320
rect 283239 336280 321560 336308
rect 283239 336277 283251 336280
rect 283193 336271 283251 336277
rect 321554 336268 321560 336280
rect 321612 336268 321618 336320
rect 348878 336268 348884 336320
rect 348936 336308 348942 336320
rect 367370 336308 367376 336320
rect 348936 336280 367376 336308
rect 348936 336268 348942 336280
rect 367370 336268 367376 336280
rect 367428 336268 367434 336320
rect 368198 336268 368204 336320
rect 368256 336308 368262 336320
rect 378781 336311 378839 336317
rect 378781 336308 378793 336311
rect 368256 336280 378793 336308
rect 368256 336268 368262 336280
rect 378781 336277 378793 336280
rect 378827 336277 378839 336311
rect 380897 336311 380955 336317
rect 380897 336308 380909 336311
rect 378781 336271 378839 336277
rect 380728 336280 380909 336308
rect 57238 336200 57244 336252
rect 57296 336240 57302 336252
rect 251266 336240 251272 336252
rect 57296 336212 251272 336240
rect 57296 336200 57302 336212
rect 251266 336200 251272 336212
rect 251324 336200 251330 336252
rect 259454 336200 259460 336252
rect 259512 336240 259518 336252
rect 261478 336240 261484 336252
rect 259512 336212 261484 336240
rect 259512 336200 259518 336212
rect 261478 336200 261484 336212
rect 261536 336200 261542 336252
rect 264882 336200 264888 336252
rect 264940 336240 264946 336252
rect 265158 336240 265164 336252
rect 264940 336212 265164 336240
rect 264940 336200 264946 336212
rect 265158 336200 265164 336212
rect 265216 336200 265222 336252
rect 269114 336200 269120 336252
rect 269172 336240 269178 336252
rect 271874 336240 271880 336252
rect 269172 336212 271880 336240
rect 269172 336200 269178 336212
rect 271874 336200 271880 336212
rect 271932 336200 271938 336252
rect 274542 336200 274548 336252
rect 274600 336240 274606 336252
rect 319254 336240 319260 336252
rect 274600 336212 319260 336240
rect 274600 336200 274606 336212
rect 319254 336200 319260 336212
rect 319312 336200 319318 336252
rect 327718 336200 327724 336252
rect 327776 336240 327782 336252
rect 328454 336240 328460 336252
rect 327776 336212 328460 336240
rect 327776 336200 327782 336212
rect 328454 336200 328460 336212
rect 328512 336200 328518 336252
rect 341610 336200 341616 336252
rect 341668 336240 341674 336252
rect 342162 336240 342168 336252
rect 341668 336212 342168 336240
rect 341668 336200 341674 336212
rect 342162 336200 342168 336212
rect 342220 336200 342226 336252
rect 346670 336200 346676 336252
rect 346728 336240 346734 336252
rect 347682 336240 347688 336252
rect 346728 336212 347688 336240
rect 346728 336200 346734 336212
rect 347682 336200 347688 336212
rect 347740 336200 347746 336252
rect 352190 336200 352196 336252
rect 352248 336240 352254 336252
rect 371786 336240 371792 336252
rect 352248 336212 371792 336240
rect 352248 336200 352254 336212
rect 371786 336200 371792 336212
rect 371844 336200 371850 336252
rect 373718 336200 373724 336252
rect 373776 336240 373782 336252
rect 374270 336240 374276 336252
rect 373776 336212 374276 336240
rect 373776 336200 373782 336212
rect 374270 336200 374276 336212
rect 374328 336200 374334 336252
rect 374380 336212 375604 336240
rect 51718 336132 51724 336184
rect 51776 336172 51782 336184
rect 247954 336172 247960 336184
rect 51776 336144 247960 336172
rect 51776 336132 51782 336144
rect 247954 336132 247960 336144
rect 248012 336132 248018 336184
rect 267642 336132 267648 336184
rect 267700 336172 267706 336184
rect 317046 336172 317052 336184
rect 267700 336144 317052 336172
rect 267700 336132 267706 336144
rect 317046 336132 317052 336144
rect 317104 336132 317110 336184
rect 351454 336132 351460 336184
rect 351512 336172 351518 336184
rect 353389 336175 353447 336181
rect 351512 336144 353340 336172
rect 351512 336132 351518 336144
rect 50338 336064 50344 336116
rect 50396 336104 50402 336116
rect 245838 336104 245844 336116
rect 50396 336076 245844 336104
rect 50396 336064 50402 336076
rect 245838 336064 245844 336076
rect 245896 336064 245902 336116
rect 270402 336064 270408 336116
rect 270460 336104 270466 336116
rect 318150 336104 318156 336116
rect 270460 336076 318156 336104
rect 270460 336064 270466 336076
rect 318150 336064 318156 336076
rect 318208 336064 318214 336116
rect 344094 336064 344100 336116
rect 344152 336104 344158 336116
rect 345658 336104 345664 336116
rect 344152 336076 345664 336104
rect 344152 336064 344158 336076
rect 345658 336064 345664 336076
rect 345716 336064 345722 336116
rect 348142 336064 348148 336116
rect 348200 336104 348206 336116
rect 349062 336104 349068 336116
rect 348200 336076 349068 336104
rect 348200 336064 348206 336076
rect 349062 336064 349068 336076
rect 349120 336064 349126 336116
rect 351086 336064 351092 336116
rect 351144 336104 351150 336116
rect 351822 336104 351828 336116
rect 351144 336076 351828 336104
rect 351144 336064 351150 336076
rect 351822 336064 351828 336076
rect 351880 336064 351886 336116
rect 352558 336064 352564 336116
rect 352616 336104 352622 336116
rect 353202 336104 353208 336116
rect 352616 336076 353208 336104
rect 352616 336064 352622 336076
rect 353202 336064 353208 336076
rect 353260 336064 353266 336116
rect 353312 336104 353340 336144
rect 353389 336141 353401 336175
rect 353435 336172 353447 336175
rect 358078 336172 358084 336184
rect 353435 336144 358084 336172
rect 353435 336141 353447 336144
rect 353389 336135 353447 336141
rect 358078 336132 358084 336144
rect 358136 336132 358142 336184
rect 363874 336132 363880 336184
rect 363932 336172 363938 336184
rect 374380 336172 374408 336212
rect 363932 336144 374408 336172
rect 363932 336132 363938 336144
rect 375466 336104 375472 336116
rect 353312 336076 375472 336104
rect 375466 336064 375472 336076
rect 375524 336064 375530 336116
rect 375576 336104 375604 336212
rect 376570 336200 376576 336252
rect 376628 336240 376634 336252
rect 380728 336240 380756 336280
rect 380897 336277 380909 336280
rect 380943 336277 380955 336311
rect 380897 336271 380955 336277
rect 381722 336268 381728 336320
rect 381780 336308 381786 336320
rect 468478 336308 468484 336320
rect 381780 336280 468484 336308
rect 381780 336268 381786 336280
rect 468478 336268 468484 336280
rect 468536 336268 468542 336320
rect 376628 336212 380756 336240
rect 376628 336200 376634 336212
rect 380802 336200 380808 336252
rect 380860 336240 380866 336252
rect 471974 336240 471980 336252
rect 380860 336212 471980 336240
rect 380860 336200 380866 336212
rect 471974 336200 471980 336212
rect 472032 336200 472038 336252
rect 378597 336175 378655 336181
rect 378597 336141 378609 336175
rect 378643 336172 378655 336175
rect 382277 336175 382335 336181
rect 382277 336172 382289 336175
rect 378643 336144 382289 336172
rect 378643 336141 378655 336144
rect 378597 336135 378655 336141
rect 382277 336141 382289 336144
rect 382323 336141 382335 336175
rect 382277 336135 382335 336141
rect 383470 336132 383476 336184
rect 383528 336172 383534 336184
rect 475378 336172 475384 336184
rect 383528 336144 475384 336172
rect 383528 336132 383534 336144
rect 475378 336132 475384 336144
rect 475436 336132 475442 336184
rect 382918 336104 382924 336116
rect 375576 336076 382924 336104
rect 382918 336064 382924 336076
rect 382976 336064 382982 336116
rect 383194 336064 383200 336116
rect 383252 336104 383258 336116
rect 478874 336104 478880 336116
rect 383252 336076 478880 336104
rect 383252 336064 383258 336076
rect 478874 336064 478880 336076
rect 478932 336064 478938 336116
rect 35158 335996 35164 336048
rect 35216 336036 35222 336048
rect 243630 336036 243636 336048
rect 35216 336008 243636 336036
rect 35216 335996 35222 336008
rect 243630 335996 243636 336008
rect 243688 335996 243694 336048
rect 263502 335996 263508 336048
rect 263560 336036 263566 336048
rect 316034 336036 316040 336048
rect 263560 336008 316040 336036
rect 263560 335996 263566 336008
rect 316034 335996 316040 336008
rect 316092 335996 316098 336048
rect 316678 335996 316684 336048
rect 316736 336036 316742 336048
rect 327258 336036 327264 336048
rect 316736 336008 327264 336036
rect 316736 335996 316742 336008
rect 327258 335996 327264 336008
rect 327316 335996 327322 336048
rect 328362 335996 328368 336048
rect 328420 336036 328426 336048
rect 335998 336036 336004 336048
rect 328420 336008 336004 336036
rect 328420 335996 328426 336008
rect 335998 335996 336004 336008
rect 336056 335996 336062 336048
rect 344830 335996 344836 336048
rect 344888 336036 344894 336048
rect 348510 336036 348516 336048
rect 344888 336008 348516 336036
rect 344888 335996 344894 336008
rect 348510 335996 348516 336008
rect 348568 335996 348574 336048
rect 353662 335996 353668 336048
rect 353720 336036 353726 336048
rect 382458 336036 382464 336048
rect 353720 336008 382464 336036
rect 353720 335996 353726 336008
rect 382458 335996 382464 336008
rect 382516 335996 382522 336048
rect 383930 335996 383936 336048
rect 383988 336036 383994 336048
rect 384850 336036 384856 336048
rect 383988 336008 384856 336036
rect 383988 335996 383994 336008
rect 384850 335996 384856 336008
rect 384908 335996 384914 336048
rect 387242 335996 387248 336048
rect 387300 336036 387306 336048
rect 387702 336036 387708 336048
rect 387300 336008 387708 336036
rect 387300 335996 387306 336008
rect 387702 335996 387708 336008
rect 387760 335996 387766 336048
rect 388346 335996 388352 336048
rect 388404 336036 388410 336048
rect 389082 336036 389088 336048
rect 388404 336008 389088 336036
rect 388404 335996 388410 336008
rect 389082 335996 389088 336008
rect 389140 335996 389146 336048
rect 389450 335996 389456 336048
rect 389508 336036 389514 336048
rect 390186 336036 390192 336048
rect 389508 336008 390192 336036
rect 389508 335996 389514 336008
rect 390186 335996 390192 336008
rect 390244 335996 390250 336048
rect 392670 335996 392676 336048
rect 392728 336036 392734 336048
rect 393130 336036 393136 336048
rect 392728 336008 393136 336036
rect 392728 335996 392734 336008
rect 393130 335996 393136 336008
rect 393188 335996 393194 336048
rect 393225 336039 393283 336045
rect 393225 336005 393237 336039
rect 393271 336036 393283 336039
rect 395338 336036 395344 336048
rect 393271 336008 395344 336036
rect 393271 336005 393283 336008
rect 393225 335999 393283 336005
rect 395338 335996 395344 336008
rect 395396 335996 395402 336048
rect 397822 335996 397828 336048
rect 397880 336036 397886 336048
rect 398558 336036 398564 336048
rect 397880 336008 398564 336036
rect 397880 335996 397886 336008
rect 398558 335996 398564 336008
rect 398616 335996 398622 336048
rect 402238 335996 402244 336048
rect 402296 336036 402302 336048
rect 402698 336036 402704 336048
rect 402296 336008 402704 336036
rect 402296 335996 402302 336008
rect 402698 335996 402704 336008
rect 402756 335996 402762 336048
rect 402793 336039 402851 336045
rect 402793 336005 402805 336039
rect 402839 336036 402851 336039
rect 497458 336036 497464 336048
rect 402839 336008 497464 336036
rect 402839 336005 402851 336008
rect 402793 335999 402851 336005
rect 497458 335996 497464 336008
rect 497516 335996 497522 336048
rect 204898 335928 204904 335980
rect 204956 335968 204962 335980
rect 276842 335968 276848 335980
rect 204956 335940 276848 335968
rect 204956 335928 204962 335940
rect 276842 335928 276848 335940
rect 276900 335928 276906 335980
rect 281350 335928 281356 335980
rect 281408 335968 281414 335980
rect 283193 335971 283251 335977
rect 283193 335968 283205 335971
rect 281408 335940 283205 335968
rect 281408 335928 281414 335940
rect 283193 335937 283205 335940
rect 283239 335937 283251 335971
rect 283193 335931 283251 335937
rect 286410 335928 286416 335980
rect 286468 335968 286474 335980
rect 315206 335968 315212 335980
rect 286468 335940 315212 335968
rect 286468 335928 286474 335940
rect 315206 335928 315212 335940
rect 315264 335928 315270 335980
rect 346302 335928 346308 335980
rect 346360 335968 346366 335980
rect 347130 335968 347136 335980
rect 346360 335940 347136 335968
rect 346360 335928 346366 335940
rect 347130 335928 347136 335940
rect 347188 335928 347194 335980
rect 356882 335928 356888 335980
rect 356940 335968 356946 335980
rect 357342 335968 357348 335980
rect 356940 335940 357348 335968
rect 356940 335928 356946 335940
rect 357342 335928 357348 335940
rect 357400 335928 357406 335980
rect 369302 335928 369308 335980
rect 369360 335968 369366 335980
rect 432598 335968 432604 335980
rect 369360 335940 432604 335968
rect 369360 335928 369366 335940
rect 432598 335928 432604 335940
rect 432656 335928 432662 335980
rect 224218 335860 224224 335912
rect 224276 335900 224282 335912
rect 291194 335900 291200 335912
rect 224276 335872 291200 335900
rect 224276 335860 224282 335872
rect 291194 335860 291200 335872
rect 291252 335860 291258 335912
rect 291930 335860 291936 335912
rect 291988 335900 291994 335912
rect 311894 335900 311900 335912
rect 291988 335872 311900 335900
rect 291988 335860 291994 335872
rect 311894 335860 311900 335872
rect 311952 335860 311958 335912
rect 333238 335860 333244 335912
rect 333296 335900 333302 335912
rect 336734 335900 336740 335912
rect 333296 335872 336740 335900
rect 333296 335860 333302 335872
rect 336734 335860 336740 335872
rect 336792 335860 336798 335912
rect 364610 335860 364616 335912
rect 364668 335900 364674 335912
rect 372525 335903 372583 335909
rect 372525 335900 372537 335903
rect 364668 335872 372537 335900
rect 364668 335860 364674 335872
rect 372525 335869 372537 335872
rect 372571 335869 372583 335903
rect 372525 335863 372583 335869
rect 372982 335860 372988 335912
rect 373040 335900 373046 335912
rect 374638 335900 374644 335912
rect 373040 335872 374644 335900
rect 373040 335860 373046 335872
rect 374638 335860 374644 335872
rect 374696 335860 374702 335912
rect 378689 335903 378747 335909
rect 378689 335869 378701 335903
rect 378735 335900 378747 335903
rect 429194 335900 429200 335912
rect 378735 335872 429200 335900
rect 378735 335869 378747 335872
rect 378689 335863 378747 335869
rect 429194 335860 429200 335872
rect 429252 335860 429258 335912
rect 233878 335792 233884 335844
rect 233936 335832 233942 335844
rect 300210 335832 300216 335844
rect 233936 335804 300216 335832
rect 233936 335792 233942 335804
rect 300210 335792 300216 335804
rect 300268 335792 300274 335844
rect 335998 335792 336004 335844
rect 336056 335832 336062 335844
rect 337470 335832 337476 335844
rect 336056 335804 337476 335832
rect 336056 335792 336062 335804
rect 337470 335792 337476 335804
rect 337528 335792 337534 335844
rect 361022 335792 361028 335844
rect 361080 335832 361086 335844
rect 361482 335832 361488 335844
rect 361080 335804 361488 335832
rect 361080 335792 361086 335804
rect 361482 335792 361488 335804
rect 361540 335792 361546 335844
rect 366450 335792 366456 335844
rect 366508 335832 366514 335844
rect 367002 335832 367008 335844
rect 366508 335804 367008 335832
rect 366508 335792 366514 335804
rect 367002 335792 367008 335804
rect 367060 335792 367066 335844
rect 367462 335792 367468 335844
rect 367520 335832 367526 335844
rect 368290 335832 368296 335844
rect 367520 335804 368296 335832
rect 367520 335792 367526 335804
rect 368290 335792 368296 335804
rect 368348 335792 368354 335844
rect 378781 335835 378839 335841
rect 378781 335801 378793 335835
rect 378827 335832 378839 335835
rect 428458 335832 428464 335844
rect 378827 335804 428464 335832
rect 378827 335801 378839 335804
rect 378781 335795 378839 335801
rect 428458 335792 428464 335804
rect 428516 335792 428522 335844
rect 222838 335724 222844 335776
rect 222896 335764 222902 335776
rect 287790 335764 287796 335776
rect 222896 335736 287796 335764
rect 222896 335724 222902 335736
rect 287790 335724 287796 335736
rect 287848 335724 287854 335776
rect 289078 335724 289084 335776
rect 289136 335764 289142 335776
rect 312998 335764 313004 335776
rect 289136 335736 313004 335764
rect 289136 335724 289142 335736
rect 312998 335724 313004 335736
rect 313056 335724 313062 335776
rect 366818 335724 366824 335776
rect 366876 335764 366882 335776
rect 425054 335764 425060 335776
rect 366876 335736 425060 335764
rect 366876 335724 366882 335736
rect 425054 335724 425060 335736
rect 425112 335724 425118 335776
rect 213178 335656 213184 335708
rect 213236 335696 213242 335708
rect 273898 335696 273904 335708
rect 213236 335668 273904 335696
rect 213236 335656 213242 335668
rect 273898 335656 273904 335668
rect 273956 335656 273962 335708
rect 288342 335656 288348 335708
rect 288400 335696 288406 335708
rect 294509 335699 294567 335705
rect 294509 335696 294521 335699
rect 288400 335668 294521 335696
rect 288400 335656 288406 335668
rect 294509 335665 294521 335668
rect 294555 335665 294567 335699
rect 294509 335659 294567 335665
rect 295978 335656 295984 335708
rect 296036 335696 296042 335708
rect 296036 335668 306374 335696
rect 296036 335656 296042 335668
rect 228358 335588 228364 335640
rect 228416 335628 228422 335640
rect 288894 335628 288900 335640
rect 228416 335600 288900 335628
rect 228416 335588 228422 335600
rect 288894 335588 288900 335600
rect 288952 335588 288958 335640
rect 296438 335588 296444 335640
rect 296496 335628 296502 335640
rect 298094 335628 298100 335640
rect 296496 335600 298100 335628
rect 296496 335588 296502 335600
rect 298094 335588 298100 335600
rect 298152 335588 298158 335640
rect 306346 335628 306374 335668
rect 310514 335656 310520 335708
rect 310572 335696 310578 335708
rect 310790 335696 310796 335708
rect 310572 335668 310796 335696
rect 310572 335656 310578 335668
rect 310790 335656 310796 335668
rect 310848 335656 310854 335708
rect 360562 335656 360568 335708
rect 360620 335696 360626 335708
rect 361298 335696 361304 335708
rect 360620 335668 361304 335696
rect 360620 335656 360626 335668
rect 361298 335656 361304 335668
rect 361356 335656 361362 335708
rect 368934 335656 368940 335708
rect 368992 335696 368998 335708
rect 369762 335696 369768 335708
rect 368992 335668 369768 335696
rect 368992 335656 368998 335668
rect 369762 335656 369768 335668
rect 369820 335656 369826 335708
rect 413097 335699 413155 335705
rect 413097 335696 413109 335699
rect 369964 335668 413109 335696
rect 314930 335628 314936 335640
rect 306346 335600 314936 335628
rect 314930 335588 314936 335600
rect 314988 335588 314994 335640
rect 366082 335588 366088 335640
rect 366140 335628 366146 335640
rect 369964 335628 369992 335668
rect 413097 335665 413109 335668
rect 413143 335665 413155 335699
rect 413097 335659 413155 335665
rect 413186 335656 413192 335708
rect 413244 335696 413250 335708
rect 413830 335696 413836 335708
rect 413244 335668 413836 335696
rect 413244 335656 413250 335668
rect 413830 335656 413836 335668
rect 413888 335656 413894 335708
rect 414750 335656 414756 335708
rect 414808 335696 414814 335708
rect 415302 335696 415308 335708
rect 414808 335668 415308 335696
rect 414808 335656 414814 335668
rect 415302 335656 415308 335668
rect 415360 335656 415366 335708
rect 372525 335631 372583 335637
rect 366140 335600 369992 335628
rect 371804 335600 372476 335628
rect 366140 335588 366146 335600
rect 231118 335520 231124 335572
rect 231176 335560 231182 335572
rect 285674 335560 285680 335572
rect 231176 335532 285680 335560
rect 231176 335520 231182 335532
rect 285674 335520 285680 335532
rect 285732 335520 285738 335572
rect 344462 335520 344468 335572
rect 344520 335560 344526 335572
rect 346946 335560 346952 335572
rect 344520 335532 346952 335560
rect 344520 335520 344526 335532
rect 346946 335520 346952 335532
rect 347004 335520 347010 335572
rect 352926 335520 352932 335572
rect 352984 335560 352990 335572
rect 353110 335560 353116 335572
rect 352984 335532 353116 335560
rect 352984 335520 352990 335532
rect 353110 335520 353116 335532
rect 353168 335520 353174 335572
rect 364978 335520 364984 335572
rect 365036 335560 365042 335572
rect 371804 335560 371832 335600
rect 365036 335532 371832 335560
rect 365036 335520 365042 335532
rect 371878 335520 371884 335572
rect 371936 335560 371942 335572
rect 372338 335560 372344 335572
rect 371936 335532 372344 335560
rect 371936 335520 371942 335532
rect 372338 335520 372344 335532
rect 372396 335520 372402 335572
rect 372448 335560 372476 335600
rect 372525 335597 372537 335631
rect 372571 335628 372583 335631
rect 414569 335631 414627 335637
rect 414569 335628 414581 335631
rect 372571 335600 414581 335628
rect 372571 335597 372583 335600
rect 372525 335591 372583 335597
rect 414569 335597 414581 335600
rect 414615 335597 414627 335631
rect 414569 335591 414627 335597
rect 414658 335588 414664 335640
rect 414716 335628 414722 335640
rect 415210 335628 415216 335640
rect 414716 335600 415216 335628
rect 414716 335588 414722 335600
rect 415210 335588 415216 335600
rect 415268 335588 415274 335640
rect 417510 335560 417516 335572
rect 372448 335532 417516 335560
rect 417510 335520 417516 335532
rect 417568 335520 417574 335572
rect 232498 335452 232504 335504
rect 232556 335492 232562 335504
rect 282362 335492 282368 335504
rect 232556 335464 282368 335492
rect 232556 335452 232562 335464
rect 282362 335452 282368 335464
rect 282420 335452 282426 335504
rect 366910 335452 366916 335504
rect 366968 335492 366974 335504
rect 418798 335492 418804 335504
rect 366968 335464 418804 335492
rect 366968 335452 366974 335464
rect 418798 335452 418804 335464
rect 418856 335452 418862 335504
rect 233970 335384 233976 335436
rect 234028 335424 234034 335436
rect 273530 335424 273536 335436
rect 234028 335396 273536 335424
rect 234028 335384 234034 335396
rect 273530 335384 273536 335396
rect 273588 335384 273594 335436
rect 341978 335384 341984 335436
rect 342036 335424 342042 335436
rect 345198 335424 345204 335436
rect 342036 335396 345204 335424
rect 342036 335384 342042 335396
rect 345198 335384 345204 335396
rect 345256 335384 345262 335436
rect 350074 335384 350080 335436
rect 350132 335424 350138 335436
rect 350350 335424 350356 335436
rect 350132 335396 350356 335424
rect 350132 335384 350138 335396
rect 350350 335384 350356 335396
rect 350408 335384 350414 335436
rect 357434 335384 357440 335436
rect 357492 335424 357498 335436
rect 393133 335427 393191 335433
rect 393133 335424 393145 335427
rect 357492 335396 393145 335424
rect 357492 335384 357498 335396
rect 393133 335393 393145 335396
rect 393179 335393 393191 335427
rect 393133 335387 393191 335393
rect 401870 335384 401876 335436
rect 401928 335424 401934 335436
rect 402606 335424 402612 335436
rect 401928 335396 402612 335424
rect 401928 335384 401934 335396
rect 402606 335384 402612 335396
rect 402664 335384 402670 335436
rect 403986 335384 403992 335436
rect 404044 335424 404050 335436
rect 404262 335424 404268 335436
rect 404044 335396 404268 335424
rect 404044 335384 404050 335396
rect 404262 335384 404268 335396
rect 404320 335384 404326 335436
rect 404722 335384 404728 335436
rect 404780 335424 404786 335436
rect 405274 335424 405280 335436
rect 404780 335396 405280 335424
rect 404780 335384 404786 335396
rect 405274 335384 405280 335396
rect 405332 335384 405338 335436
rect 405366 335384 405372 335436
rect 405424 335424 405430 335436
rect 405550 335424 405556 335436
rect 405424 335396 405556 335424
rect 405424 335384 405430 335396
rect 405550 335384 405556 335396
rect 405608 335384 405614 335436
rect 406562 335384 406568 335436
rect 406620 335424 406626 335436
rect 406838 335424 406844 335436
rect 406620 335396 406844 335424
rect 406620 335384 406626 335396
rect 406838 335384 406844 335396
rect 406896 335384 406902 335436
rect 407666 335384 407672 335436
rect 407724 335424 407730 335436
rect 408310 335424 408316 335436
rect 407724 335396 408316 335424
rect 407724 335384 407730 335396
rect 408310 335384 408316 335396
rect 408368 335384 408374 335436
rect 409506 335384 409512 335436
rect 409564 335424 409570 335436
rect 409782 335424 409788 335436
rect 409564 335396 409788 335424
rect 409564 335384 409570 335396
rect 409782 335384 409788 335396
rect 409840 335384 409846 335436
rect 410702 335384 410708 335436
rect 410760 335424 410766 335436
rect 411070 335424 411076 335436
rect 410760 335396 411076 335424
rect 410760 335384 410766 335396
rect 411070 335384 411076 335396
rect 411128 335384 411134 335436
rect 412082 335384 412088 335436
rect 412140 335424 412146 335436
rect 412358 335424 412364 335436
rect 412140 335396 412364 335424
rect 412140 335384 412146 335396
rect 412358 335384 412364 335396
rect 412416 335384 412422 335436
rect 414569 335427 414627 335433
rect 414569 335393 414581 335427
rect 414615 335424 414627 335427
rect 418154 335424 418160 335436
rect 414615 335396 418160 335424
rect 414615 335393 414627 335396
rect 414569 335387 414627 335393
rect 418154 335384 418160 335396
rect 418212 335384 418218 335436
rect 274450 335316 274456 335368
rect 274508 335356 274514 335368
rect 278774 335356 278780 335368
rect 274508 335328 278780 335356
rect 274508 335316 274514 335328
rect 278774 335316 278780 335328
rect 278832 335316 278838 335368
rect 289998 335356 290004 335368
rect 289786 335328 290004 335356
rect 179322 335248 179328 335300
rect 179380 335288 179386 335300
rect 289786 335288 289814 335328
rect 289998 335316 290004 335328
rect 290056 335316 290062 335368
rect 332502 335316 332508 335368
rect 332560 335356 332566 335368
rect 337102 335356 337108 335368
rect 332560 335328 337108 335356
rect 332560 335316 332566 335328
rect 337102 335316 337108 335328
rect 337160 335316 337166 335368
rect 344922 335316 344928 335368
rect 344980 335356 344986 335368
rect 345750 335356 345756 335368
rect 344980 335328 345756 335356
rect 344980 335316 344986 335328
rect 345750 335316 345756 335328
rect 345808 335316 345814 335368
rect 355410 335316 355416 335368
rect 355468 335356 355474 335368
rect 388438 335356 388444 335368
rect 355468 335328 388444 335356
rect 355468 335316 355474 335328
rect 388438 335316 388444 335328
rect 388496 335316 388502 335368
rect 388806 335316 388812 335368
rect 388864 335356 388870 335368
rect 402793 335359 402851 335365
rect 402793 335356 402805 335359
rect 388864 335328 402805 335356
rect 388864 335316 388870 335328
rect 402793 335325 402805 335328
rect 402839 335325 402851 335359
rect 402793 335319 402851 335325
rect 403250 335316 403256 335368
rect 403308 335356 403314 335368
rect 404170 335356 404176 335368
rect 403308 335328 404176 335356
rect 403308 335316 403314 335328
rect 404170 335316 404176 335328
rect 404228 335316 404234 335368
rect 405090 335316 405096 335368
rect 405148 335356 405154 335368
rect 405642 335356 405648 335368
rect 405148 335328 405648 335356
rect 405148 335316 405154 335328
rect 405642 335316 405648 335328
rect 405700 335316 405706 335368
rect 406194 335316 406200 335368
rect 406252 335356 406258 335368
rect 407022 335356 407028 335368
rect 406252 335328 407028 335356
rect 406252 335316 406258 335328
rect 407022 335316 407028 335328
rect 407080 335316 407086 335368
rect 408770 335316 408776 335368
rect 408828 335356 408834 335368
rect 409598 335356 409604 335368
rect 408828 335328 409604 335356
rect 408828 335316 408834 335328
rect 409598 335316 409604 335328
rect 409656 335316 409662 335368
rect 410242 335316 410248 335368
rect 410300 335356 410306 335368
rect 410978 335356 410984 335368
rect 410300 335328 410984 335356
rect 410300 335316 410306 335328
rect 410978 335316 410984 335328
rect 411036 335316 411042 335368
rect 411714 335316 411720 335368
rect 411772 335356 411778 335368
rect 412450 335356 412456 335368
rect 411772 335328 412456 335356
rect 411772 335316 411778 335328
rect 412450 335316 412456 335328
rect 412508 335316 412514 335368
rect 413097 335359 413155 335365
rect 413097 335325 413109 335359
rect 413143 335356 413155 335359
rect 421558 335356 421564 335368
rect 413143 335328 421564 335356
rect 413143 335325 413155 335328
rect 413097 335319 413155 335325
rect 421558 335316 421564 335328
rect 421616 335316 421622 335368
rect 179380 335260 289814 335288
rect 179380 335248 179386 335260
rect 388990 335248 388996 335300
rect 389048 335288 389054 335300
rect 483014 335288 483020 335300
rect 389048 335260 483020 335288
rect 389048 335248 389054 335260
rect 483014 335248 483020 335260
rect 483072 335248 483078 335300
rect 169662 335180 169668 335232
rect 169720 335220 169726 335232
rect 286686 335220 286692 335232
rect 169720 335192 286692 335220
rect 169720 335180 169726 335192
rect 286686 335180 286692 335192
rect 286744 335180 286750 335232
rect 384298 335180 384304 335232
rect 384356 335220 384362 335232
rect 481634 335220 481640 335232
rect 384356 335192 481640 335220
rect 384356 335180 384362 335192
rect 481634 335180 481640 335192
rect 481692 335180 481698 335232
rect 161382 335112 161388 335164
rect 161440 335152 161446 335164
rect 284478 335152 284484 335164
rect 161440 335124 284484 335152
rect 161440 335112 161446 335124
rect 284478 335112 284484 335124
rect 284536 335112 284542 335164
rect 391934 335112 391940 335164
rect 391992 335152 391998 335164
rect 490006 335152 490012 335164
rect 391992 335124 490012 335152
rect 391992 335112 391998 335124
rect 490006 335112 490012 335124
rect 490064 335112 490070 335164
rect 144822 335044 144828 335096
rect 144880 335084 144886 335096
rect 276014 335084 276020 335096
rect 144880 335056 276020 335084
rect 144880 335044 144886 335056
rect 276014 335044 276020 335056
rect 276072 335044 276078 335096
rect 390094 335044 390100 335096
rect 390152 335084 390158 335096
rect 500954 335084 500960 335096
rect 390152 335056 500960 335084
rect 390152 335044 390158 335056
rect 500954 335044 500960 335056
rect 501012 335044 501018 335096
rect 147582 334976 147588 335028
rect 147640 335016 147646 335028
rect 280246 335016 280252 335028
rect 147640 334988 280252 335016
rect 147640 334976 147646 334988
rect 280246 334976 280252 334988
rect 280304 334976 280310 335028
rect 392302 334976 392308 335028
rect 392360 335016 392366 335028
rect 507854 335016 507860 335028
rect 392360 334988 507860 335016
rect 392360 334976 392366 334988
rect 507854 334976 507860 334988
rect 507912 334976 507918 335028
rect 140682 334908 140688 334960
rect 140740 334948 140746 334960
rect 277946 334948 277952 334960
rect 140740 334920 277952 334948
rect 140740 334908 140746 334920
rect 277946 334908 277952 334920
rect 278004 334908 278010 334960
rect 393774 334908 393780 334960
rect 393832 334948 393838 334960
rect 512638 334948 512644 334960
rect 393832 334920 512644 334948
rect 393832 334908 393838 334920
rect 512638 334908 512644 334920
rect 512696 334908 512702 334960
rect 86862 334840 86868 334892
rect 86920 334880 86926 334892
rect 259454 334880 259460 334892
rect 86920 334852 259460 334880
rect 86920 334840 86926 334852
rect 259454 334840 259460 334852
rect 259512 334840 259518 334892
rect 395890 334840 395896 334892
rect 395948 334880 395954 334892
rect 520274 334880 520280 334892
rect 395948 334852 520280 334880
rect 395948 334840 395954 334852
rect 520274 334840 520280 334852
rect 520332 334840 520338 334892
rect 87598 334772 87604 334824
rect 87656 334812 87662 334824
rect 260926 334812 260932 334824
rect 87656 334784 260932 334812
rect 87656 334772 87662 334784
rect 260926 334772 260932 334784
rect 260984 334772 260990 334824
rect 398190 334772 398196 334824
rect 398248 334812 398254 334824
rect 526438 334812 526444 334824
rect 398248 334784 526444 334812
rect 398248 334772 398254 334784
rect 526438 334772 526444 334784
rect 526496 334772 526502 334824
rect 54478 334704 54484 334756
rect 54536 334744 54542 334756
rect 247586 334744 247592 334756
rect 54536 334716 247592 334744
rect 54536 334704 54542 334716
rect 247586 334704 247592 334716
rect 247644 334704 247650 334756
rect 397086 334704 397092 334756
rect 397144 334744 397150 334756
rect 522298 334744 522304 334756
rect 397144 334716 522304 334744
rect 397144 334704 397150 334716
rect 522298 334704 522304 334716
rect 522356 334704 522362 334756
rect 29638 334636 29644 334688
rect 29696 334676 29702 334688
rect 243262 334676 243268 334688
rect 29696 334648 243268 334676
rect 29696 334636 29702 334648
rect 243262 334636 243268 334648
rect 243320 334636 243326 334688
rect 398466 334636 398472 334688
rect 398524 334676 398530 334688
rect 528554 334676 528560 334688
rect 398524 334648 528560 334676
rect 398524 334636 398530 334648
rect 528554 334636 528560 334648
rect 528612 334636 528618 334688
rect 22738 334568 22744 334620
rect 22796 334608 22802 334620
rect 238846 334608 238852 334620
rect 22796 334580 238852 334608
rect 22796 334568 22802 334580
rect 238846 334568 238852 334580
rect 238904 334568 238910 334620
rect 402514 334568 402520 334620
rect 402572 334608 402578 334620
rect 540238 334608 540244 334620
rect 402572 334580 540244 334608
rect 402572 334568 402578 334580
rect 540238 334568 540244 334580
rect 540296 334568 540302 334620
rect 197262 334500 197268 334552
rect 197320 334540 197326 334552
rect 292482 334540 292488 334552
rect 197320 334512 292488 334540
rect 197320 334500 197326 334512
rect 292482 334500 292488 334512
rect 292540 334500 292546 334552
rect 374270 334500 374276 334552
rect 374328 334540 374334 334552
rect 448514 334540 448520 334552
rect 374328 334512 448520 334540
rect 374328 334500 374334 334512
rect 448514 334500 448520 334512
rect 448572 334500 448578 334552
rect 202782 334432 202788 334484
rect 202840 334472 202846 334484
rect 296530 334472 296536 334484
rect 202840 334444 296536 334472
rect 202840 334432 202846 334444
rect 296530 334432 296536 334444
rect 296588 334432 296594 334484
rect 371510 334432 371516 334484
rect 371568 334472 371574 334484
rect 440326 334472 440332 334484
rect 371568 334444 440332 334472
rect 371568 334432 371574 334444
rect 440326 334432 440332 334444
rect 440384 334432 440390 334484
rect 216582 334364 216588 334416
rect 216640 334404 216646 334416
rect 300486 334404 300492 334416
rect 216640 334376 300492 334404
rect 216640 334364 216646 334376
rect 300486 334364 300492 334376
rect 300544 334364 300550 334416
rect 223482 334296 223488 334348
rect 223540 334336 223546 334348
rect 303614 334336 303620 334348
rect 223540 334308 303620 334336
rect 223540 334296 223546 334308
rect 303614 334296 303620 334308
rect 303672 334296 303678 334348
rect 205542 333888 205548 333940
rect 205600 333928 205606 333940
rect 296438 333928 296444 333940
rect 205600 333900 296444 333928
rect 205600 333888 205606 333900
rect 296438 333888 296444 333900
rect 296496 333888 296502 333940
rect 374638 333888 374644 333940
rect 374696 333928 374702 333940
rect 445754 333928 445760 333940
rect 374696 333900 445760 333928
rect 374696 333888 374702 333900
rect 445754 333888 445760 333900
rect 445812 333888 445818 333940
rect 198642 333820 198648 333872
rect 198700 333860 198706 333872
rect 295794 333860 295800 333872
rect 198700 333832 295800 333860
rect 198700 333820 198706 333832
rect 295794 333820 295800 333832
rect 295852 333820 295858 333872
rect 373810 333820 373816 333872
rect 373868 333860 373874 333872
rect 448606 333860 448612 333872
rect 373868 333832 448612 333860
rect 373868 333820 373874 333832
rect 448606 333820 448612 333832
rect 448664 333820 448670 333872
rect 177942 333752 177948 333804
rect 178000 333792 178006 333804
rect 288434 333792 288440 333804
rect 178000 333764 288440 333792
rect 178000 333752 178006 333764
rect 288434 333752 288440 333764
rect 288492 333752 288498 333804
rect 375006 333752 375012 333804
rect 375064 333792 375070 333804
rect 452654 333792 452660 333804
rect 375064 333764 452660 333792
rect 375064 333752 375070 333764
rect 452654 333752 452660 333764
rect 452712 333752 452718 333804
rect 162762 333684 162768 333736
rect 162820 333724 162826 333736
rect 284846 333724 284852 333736
rect 162820 333696 284852 333724
rect 162820 333684 162826 333696
rect 284846 333684 284852 333696
rect 284904 333684 284910 333736
rect 377398 333684 377404 333736
rect 377456 333724 377462 333736
rect 459554 333724 459560 333736
rect 377456 333696 459560 333724
rect 377456 333684 377462 333696
rect 459554 333684 459560 333696
rect 459612 333684 459618 333736
rect 158622 333616 158628 333668
rect 158680 333656 158686 333668
rect 282638 333656 282644 333668
rect 158680 333628 282644 333656
rect 158680 333616 158686 333628
rect 282638 333616 282644 333628
rect 282696 333616 282702 333668
rect 380526 333616 380532 333668
rect 380584 333656 380590 333668
rect 470594 333656 470600 333668
rect 380584 333628 470600 333656
rect 380584 333616 380590 333628
rect 470594 333616 470600 333628
rect 470652 333616 470658 333668
rect 151722 333548 151728 333600
rect 151780 333588 151786 333600
rect 281442 333588 281448 333600
rect 151780 333560 281448 333588
rect 151780 333548 151786 333560
rect 281442 333548 281448 333560
rect 281500 333548 281506 333600
rect 387610 333548 387616 333600
rect 387668 333588 387674 333600
rect 492674 333588 492680 333600
rect 387668 333560 492680 333588
rect 387668 333548 387674 333560
rect 492674 333548 492680 333560
rect 492732 333548 492738 333600
rect 104158 333480 104164 333532
rect 104216 333520 104222 333532
rect 266354 333520 266360 333532
rect 104216 333492 266360 333520
rect 104216 333480 104222 333492
rect 266354 333480 266360 333492
rect 266412 333480 266418 333532
rect 390922 333480 390928 333532
rect 390980 333520 390986 333532
rect 502978 333520 502984 333532
rect 390980 333492 502984 333520
rect 390980 333480 390986 333492
rect 502978 333480 502984 333492
rect 503036 333480 503042 333532
rect 93118 333412 93124 333464
rect 93176 333452 93182 333464
rect 262950 333452 262956 333464
rect 93176 333424 262956 333452
rect 93176 333412 93182 333424
rect 262950 333412 262956 333424
rect 263008 333412 263014 333464
rect 394602 333412 394608 333464
rect 394660 333452 394666 333464
rect 515398 333452 515404 333464
rect 394660 333424 515404 333452
rect 394660 333412 394666 333424
rect 515398 333412 515404 333424
rect 515456 333412 515462 333464
rect 88978 333344 88984 333396
rect 89036 333384 89042 333396
rect 261938 333384 261944 333396
rect 89036 333356 261944 333384
rect 89036 333344 89042 333356
rect 261938 333344 261944 333356
rect 261996 333344 262002 333396
rect 399294 333344 399300 333396
rect 399352 333384 399358 333396
rect 530578 333384 530584 333396
rect 399352 333356 530584 333384
rect 399352 333344 399358 333356
rect 530578 333344 530584 333356
rect 530636 333344 530642 333396
rect 84102 333276 84108 333328
rect 84160 333316 84166 333328
rect 251269 333319 251327 333325
rect 251269 333316 251281 333319
rect 84160 333288 251281 333316
rect 84160 333276 84166 333288
rect 251269 333285 251281 333288
rect 251315 333285 251327 333319
rect 251269 333279 251327 333285
rect 400122 333276 400128 333328
rect 400180 333316 400186 333328
rect 533338 333316 533344 333328
rect 400180 333288 533344 333316
rect 400180 333276 400186 333288
rect 533338 333276 533344 333288
rect 533396 333276 533402 333328
rect 39298 333208 39304 333260
rect 39356 333248 39362 333260
rect 241790 333248 241796 333260
rect 39356 333220 241796 333248
rect 39356 333208 39362 333220
rect 241790 333208 241796 333220
rect 241848 333208 241854 333260
rect 401502 333208 401508 333260
rect 401560 333248 401566 333260
rect 538214 333248 538220 333260
rect 401560 333220 538220 333248
rect 401560 333208 401566 333220
rect 538214 333208 538220 333220
rect 538272 333208 538278 333260
rect 209682 333140 209688 333192
rect 209740 333180 209746 333192
rect 299106 333180 299112 333192
rect 209740 333152 299112 333180
rect 209740 333140 209746 333152
rect 299106 333140 299112 333152
rect 299164 333140 299170 333192
rect 227622 333072 227628 333124
rect 227680 333112 227686 333124
rect 304626 333112 304632 333124
rect 227680 333084 304632 333112
rect 227680 333072 227686 333084
rect 304626 333072 304632 333084
rect 304684 333072 304690 333124
rect 251269 333047 251327 333053
rect 251269 333013 251281 333047
rect 251315 333044 251327 333047
rect 260374 333044 260380 333056
rect 251315 333016 260380 333044
rect 251315 333013 251327 333016
rect 251269 333007 251327 333013
rect 260374 333004 260380 333016
rect 260432 333004 260438 333056
rect 219250 332528 219256 332580
rect 219308 332568 219314 332580
rect 302602 332568 302608 332580
rect 219308 332540 302608 332568
rect 219308 332528 219314 332540
rect 302602 332528 302608 332540
rect 302660 332528 302666 332580
rect 188982 332460 188988 332512
rect 189040 332500 189046 332512
rect 291562 332500 291568 332512
rect 189040 332472 291568 332500
rect 189040 332460 189046 332472
rect 291562 332460 291568 332472
rect 291620 332460 291626 332512
rect 182082 332392 182088 332444
rect 182140 332432 182146 332444
rect 290826 332432 290832 332444
rect 182140 332404 290832 332432
rect 182140 332392 182146 332404
rect 290826 332392 290832 332404
rect 290884 332392 290890 332444
rect 175182 332324 175188 332376
rect 175240 332364 175246 332376
rect 288526 332364 288532 332376
rect 175240 332336 288532 332364
rect 175240 332324 175246 332336
rect 288526 332324 288532 332336
rect 288584 332324 288590 332376
rect 376202 332324 376208 332376
rect 376260 332364 376266 332376
rect 456886 332364 456892 332376
rect 376260 332336 456892 332364
rect 376260 332324 376266 332336
rect 456886 332324 456892 332336
rect 456944 332324 456950 332376
rect 171042 332256 171048 332308
rect 171100 332296 171106 332308
rect 287422 332296 287428 332308
rect 171100 332268 287428 332296
rect 171100 332256 171106 332268
rect 287422 332256 287428 332268
rect 287480 332256 287486 332308
rect 378502 332256 378508 332308
rect 378560 332296 378566 332308
rect 463694 332296 463700 332308
rect 378560 332268 463700 332296
rect 378560 332256 378566 332268
rect 463694 332256 463700 332268
rect 463752 332256 463758 332308
rect 143442 332188 143448 332240
rect 143500 332228 143506 332240
rect 274450 332228 274456 332240
rect 143500 332200 274456 332228
rect 143500 332188 143506 332200
rect 274450 332188 274456 332200
rect 274508 332188 274514 332240
rect 379422 332188 379428 332240
rect 379480 332228 379486 332240
rect 466454 332228 466460 332240
rect 379480 332200 466460 332228
rect 379480 332188 379486 332200
rect 466454 332188 466460 332200
rect 466512 332188 466518 332240
rect 124122 332120 124128 332172
rect 124180 332160 124186 332172
rect 271782 332160 271788 332172
rect 124180 332132 271788 332160
rect 124180 332120 124186 332132
rect 271782 332120 271788 332132
rect 271840 332120 271846 332172
rect 382826 332120 382832 332172
rect 382884 332160 382890 332172
rect 477494 332160 477500 332172
rect 382884 332132 477500 332160
rect 382884 332120 382890 332132
rect 477494 332120 477500 332132
rect 477552 332120 477558 332172
rect 106182 332052 106188 332104
rect 106240 332092 106246 332104
rect 267366 332092 267372 332104
rect 106240 332064 267372 332092
rect 106240 332052 106246 332064
rect 267366 332052 267372 332064
rect 267424 332052 267430 332104
rect 385310 332052 385316 332104
rect 385368 332092 385374 332104
rect 485774 332092 485780 332104
rect 385368 332064 485780 332092
rect 385368 332052 385374 332064
rect 485774 332052 485780 332064
rect 485832 332052 485838 332104
rect 99282 331984 99288 332036
rect 99340 332024 99346 332036
rect 264882 332024 264888 332036
rect 99340 331996 264888 332024
rect 99340 331984 99346 331996
rect 264882 331984 264888 331996
rect 264940 331984 264946 332036
rect 386322 331984 386328 332036
rect 386380 332024 386386 332036
rect 489178 332024 489184 332036
rect 386380 331996 489184 332024
rect 386380 331984 386386 331996
rect 489178 331984 489184 331996
rect 489236 331984 489242 332036
rect 95142 331916 95148 331968
rect 95200 331956 95206 331968
rect 264054 331956 264060 331968
rect 95200 331928 264060 331956
rect 95200 331916 95206 331928
rect 264054 331916 264060 331928
rect 264112 331916 264118 331968
rect 388714 331916 388720 331968
rect 388772 331956 388778 331968
rect 496814 331956 496820 331968
rect 388772 331928 496820 331956
rect 388772 331916 388778 331928
rect 496814 331916 496820 331928
rect 496872 331916 496878 331968
rect 68278 331848 68284 331900
rect 68336 331888 68342 331900
rect 250162 331888 250168 331900
rect 68336 331860 250168 331888
rect 68336 331848 68342 331860
rect 250162 331848 250168 331860
rect 250220 331848 250226 331900
rect 391842 331848 391848 331900
rect 391900 331888 391906 331900
rect 506474 331888 506480 331900
rect 391900 331860 506480 331888
rect 391900 331848 391906 331860
rect 506474 331848 506480 331860
rect 506532 331848 506538 331900
rect 410610 331100 410616 331152
rect 410668 331140 410674 331152
rect 411162 331140 411168 331152
rect 410668 331112 411168 331140
rect 410668 331100 410674 331112
rect 411162 331100 411168 331112
rect 411220 331100 411226 331152
rect 153102 330964 153108 331016
rect 153160 331004 153166 331016
rect 281994 331004 282000 331016
rect 153160 330976 282000 331004
rect 153160 330964 153166 330976
rect 281994 330964 282000 330976
rect 282052 330964 282058 331016
rect 146202 330896 146208 330948
rect 146260 330936 146266 330948
rect 277854 330936 277860 330948
rect 146260 330908 277860 330936
rect 146260 330896 146266 330908
rect 277854 330896 277860 330908
rect 277912 330896 277918 330948
rect 117222 330828 117228 330880
rect 117280 330868 117286 330880
rect 270862 330868 270868 330880
rect 117280 330840 270868 330868
rect 117280 330828 117286 330840
rect 270862 330828 270868 330840
rect 270920 330828 270926 330880
rect 399662 330828 399668 330880
rect 399720 330868 399726 330880
rect 485038 330868 485044 330880
rect 399720 330840 485044 330868
rect 399720 330828 399726 330840
rect 485038 330828 485044 330840
rect 485096 330828 485102 330880
rect 113082 330760 113088 330812
rect 113140 330800 113146 330812
rect 269574 330800 269580 330812
rect 113140 330772 269580 330800
rect 113140 330760 113146 330772
rect 269574 330760 269580 330772
rect 269632 330760 269638 330812
rect 331582 330760 331588 330812
rect 331640 330760 331646 330812
rect 389818 330760 389824 330812
rect 389876 330800 389882 330812
rect 499574 330800 499580 330812
rect 389876 330772 499580 330800
rect 389876 330760 389882 330772
rect 499574 330760 499580 330772
rect 499632 330760 499638 330812
rect 111058 330692 111064 330744
rect 111116 330732 111122 330744
rect 268470 330732 268476 330744
rect 111116 330704 268476 330732
rect 111116 330692 111122 330704
rect 268470 330692 268476 330704
rect 268528 330692 268534 330744
rect 81342 330624 81348 330676
rect 81400 330664 81406 330676
rect 259638 330664 259644 330676
rect 81400 330636 259644 330664
rect 81400 330624 81406 330636
rect 259638 330624 259644 330636
rect 259696 330624 259702 330676
rect 331600 330608 331628 330760
rect 392854 330692 392860 330744
rect 392912 330732 392918 330744
rect 510614 330732 510620 330744
rect 392912 330704 510620 330732
rect 392912 330692 392918 330704
rect 510614 330692 510620 330704
rect 510672 330692 510678 330744
rect 394142 330624 394148 330676
rect 394200 330664 394206 330676
rect 514754 330664 514760 330676
rect 394200 330636 514760 330664
rect 394200 330624 394206 330636
rect 514754 330624 514760 330636
rect 514812 330624 514818 330676
rect 61378 330556 61384 330608
rect 61436 330596 61442 330608
rect 252554 330596 252560 330608
rect 61436 330568 252560 330596
rect 61436 330556 61442 330568
rect 252554 330556 252560 330568
rect 252612 330556 252618 330608
rect 331582 330556 331588 330608
rect 331640 330556 331646 330608
rect 395154 330556 395160 330608
rect 395212 330596 395218 330608
rect 517514 330596 517520 330608
rect 395212 330568 517520 330596
rect 395212 330556 395218 330568
rect 517514 330556 517520 330568
rect 517572 330556 517578 330608
rect 33778 330488 33784 330540
rect 33836 330528 33842 330540
rect 33836 330500 238754 330528
rect 33836 330488 33842 330500
rect 234798 330420 234804 330472
rect 234856 330460 234862 330472
rect 235258 330460 235264 330472
rect 234856 330432 235264 330460
rect 234856 330420 234862 330432
rect 235258 330420 235264 330432
rect 235316 330420 235322 330472
rect 236086 330420 236092 330472
rect 236144 330460 236150 330472
rect 237006 330460 237012 330472
rect 236144 330432 237012 330460
rect 236144 330420 236150 330432
rect 237006 330420 237012 330432
rect 237064 330420 237070 330472
rect 237374 330420 237380 330472
rect 237432 330460 237438 330472
rect 238478 330460 238484 330472
rect 237432 330432 238484 330460
rect 237432 330420 237438 330432
rect 238478 330420 238484 330432
rect 238536 330420 238542 330472
rect 238726 330460 238754 330500
rect 241606 330488 241612 330540
rect 241664 330528 241670 330540
rect 242526 330528 242532 330540
rect 241664 330500 242532 330528
rect 241664 330488 241670 330500
rect 242526 330488 242532 330500
rect 242584 330488 242590 330540
rect 244366 330488 244372 330540
rect 244424 330528 244430 330540
rect 245102 330528 245108 330540
rect 244424 330500 245108 330528
rect 244424 330488 244430 330500
rect 245102 330488 245108 330500
rect 245160 330488 245166 330540
rect 247126 330488 247132 330540
rect 247184 330528 247190 330540
rect 247310 330528 247316 330540
rect 247184 330500 247316 330528
rect 247184 330488 247190 330500
rect 247310 330488 247316 330500
rect 247368 330488 247374 330540
rect 248506 330488 248512 330540
rect 248564 330528 248570 330540
rect 249426 330528 249432 330540
rect 248564 330500 249432 330528
rect 248564 330488 248570 330500
rect 249426 330488 249432 330500
rect 249484 330488 249490 330540
rect 249978 330488 249984 330540
rect 250036 330528 250042 330540
rect 250898 330528 250904 330540
rect 250036 330500 250904 330528
rect 250036 330488 250042 330500
rect 250898 330488 250904 330500
rect 250956 330488 250962 330540
rect 251266 330488 251272 330540
rect 251324 330528 251330 330540
rect 252002 330528 252008 330540
rect 251324 330500 252008 330528
rect 251324 330488 251330 330500
rect 252002 330488 252008 330500
rect 252060 330488 252066 330540
rect 253934 330488 253940 330540
rect 253992 330528 253998 330540
rect 254578 330528 254584 330540
rect 253992 330500 254584 330528
rect 253992 330488 253998 330500
rect 254578 330488 254584 330500
rect 254636 330488 254642 330540
rect 255314 330488 255320 330540
rect 255372 330528 255378 330540
rect 255682 330528 255688 330540
rect 255372 330500 255688 330528
rect 255372 330488 255378 330500
rect 255682 330488 255688 330500
rect 255740 330488 255746 330540
rect 258166 330488 258172 330540
rect 258224 330528 258230 330540
rect 258994 330528 259000 330540
rect 258224 330500 259000 330528
rect 258224 330488 258230 330500
rect 258994 330488 259000 330500
rect 259052 330488 259058 330540
rect 265158 330488 265164 330540
rect 265216 330528 265222 330540
rect 265894 330528 265900 330540
rect 265216 330500 265900 330528
rect 265216 330488 265222 330500
rect 265894 330488 265900 330500
rect 265952 330488 265958 330540
rect 266446 330488 266452 330540
rect 266504 330528 266510 330540
rect 266998 330528 267004 330540
rect 266504 330500 267004 330528
rect 266504 330488 266510 330500
rect 266998 330488 267004 330500
rect 267056 330488 267062 330540
rect 270586 330488 270592 330540
rect 270644 330528 270650 330540
rect 271322 330528 271328 330540
rect 270644 330500 271328 330528
rect 270644 330488 270650 330500
rect 271322 330488 271328 330500
rect 271380 330488 271386 330540
rect 271966 330488 271972 330540
rect 272024 330528 272030 330540
rect 272426 330528 272432 330540
rect 272024 330500 272432 330528
rect 272024 330488 272030 330500
rect 272426 330488 272432 330500
rect 272484 330488 272490 330540
rect 285766 330488 285772 330540
rect 285824 330528 285830 330540
rect 286318 330528 286324 330540
rect 285824 330500 286324 330528
rect 285824 330488 285830 330500
rect 286318 330488 286324 330500
rect 286376 330488 286382 330540
rect 287146 330488 287152 330540
rect 287204 330528 287210 330540
rect 288158 330528 288164 330540
rect 287204 330500 288164 330528
rect 287204 330488 287210 330500
rect 288158 330488 288164 330500
rect 288216 330488 288222 330540
rect 291286 330488 291292 330540
rect 291344 330528 291350 330540
rect 291838 330528 291844 330540
rect 291344 330500 291844 330528
rect 291344 330488 291350 330500
rect 291838 330488 291844 330500
rect 291896 330488 291902 330540
rect 294138 330488 294144 330540
rect 294196 330528 294202 330540
rect 295150 330528 295156 330540
rect 294196 330500 295156 330528
rect 294196 330488 294202 330500
rect 295150 330488 295156 330500
rect 295208 330488 295214 330540
rect 299566 330488 299572 330540
rect 299624 330528 299630 330540
rect 300578 330528 300584 330540
rect 299624 330500 300584 330528
rect 299624 330488 299630 330500
rect 300578 330488 300584 330500
rect 300636 330488 300642 330540
rect 300946 330488 300952 330540
rect 301004 330528 301010 330540
rect 301682 330528 301688 330540
rect 301004 330500 301688 330528
rect 301004 330488 301010 330500
rect 301682 330488 301688 330500
rect 301740 330488 301746 330540
rect 311986 330488 311992 330540
rect 312044 330528 312050 330540
rect 312630 330528 312636 330540
rect 312044 330500 312636 330528
rect 312044 330488 312050 330500
rect 312630 330488 312636 330500
rect 312688 330488 312694 330540
rect 313274 330488 313280 330540
rect 313332 330528 313338 330540
rect 314102 330528 314108 330540
rect 313332 330500 314108 330528
rect 313332 330488 313338 330500
rect 314102 330488 314108 330500
rect 314160 330488 314166 330540
rect 317598 330488 317604 330540
rect 317656 330528 317662 330540
rect 318518 330528 318524 330540
rect 317656 330500 318524 330528
rect 317656 330488 317662 330500
rect 318518 330488 318524 330500
rect 318576 330488 318582 330540
rect 318886 330488 318892 330540
rect 318944 330528 318950 330540
rect 319530 330528 319536 330540
rect 318944 330500 319536 330528
rect 318944 330488 318950 330500
rect 319530 330488 319536 330500
rect 319588 330488 319594 330540
rect 320174 330488 320180 330540
rect 320232 330528 320238 330540
rect 321002 330528 321008 330540
rect 320232 330500 321008 330528
rect 320232 330488 320238 330500
rect 321002 330488 321008 330500
rect 321060 330488 321066 330540
rect 321646 330488 321652 330540
rect 321704 330528 321710 330540
rect 322106 330528 322112 330540
rect 321704 330500 322112 330528
rect 321704 330488 321710 330500
rect 322106 330488 322112 330500
rect 322164 330488 322170 330540
rect 323118 330488 323124 330540
rect 323176 330528 323182 330540
rect 323946 330528 323952 330540
rect 323176 330500 323952 330528
rect 323176 330488 323182 330500
rect 323946 330488 323952 330500
rect 324004 330488 324010 330540
rect 324314 330488 324320 330540
rect 324372 330528 324378 330540
rect 324682 330528 324688 330540
rect 324372 330500 324688 330528
rect 324372 330488 324378 330500
rect 324682 330488 324688 330500
rect 324740 330488 324746 330540
rect 325786 330488 325792 330540
rect 325844 330528 325850 330540
rect 326522 330528 326528 330540
rect 325844 330500 326528 330528
rect 325844 330488 325850 330500
rect 326522 330488 326528 330500
rect 326580 330488 326586 330540
rect 329926 330488 329932 330540
rect 329984 330528 329990 330540
rect 330938 330528 330944 330540
rect 329984 330500 330944 330528
rect 329984 330488 329990 330500
rect 330938 330488 330944 330500
rect 330996 330488 331002 330540
rect 331490 330488 331496 330540
rect 331548 330528 331554 330540
rect 331950 330528 331956 330540
rect 331548 330500 331956 330528
rect 331548 330488 331554 330500
rect 331950 330488 331956 330500
rect 332008 330488 332014 330540
rect 332594 330488 332600 330540
rect 332652 330528 332658 330540
rect 333422 330528 333428 330540
rect 332652 330500 333428 330528
rect 332652 330488 332658 330500
rect 333422 330488 333428 330500
rect 333480 330488 333486 330540
rect 334066 330488 334072 330540
rect 334124 330528 334130 330540
rect 334526 330528 334532 330540
rect 334124 330500 334532 330528
rect 334124 330488 334130 330500
rect 334526 330488 334532 330500
rect 334584 330488 334590 330540
rect 335446 330488 335452 330540
rect 335504 330528 335510 330540
rect 336366 330528 336372 330540
rect 335504 330500 336372 330528
rect 335504 330488 335510 330500
rect 336366 330488 336372 330500
rect 336424 330488 336430 330540
rect 338114 330488 338120 330540
rect 338172 330528 338178 330540
rect 338574 330528 338580 330540
rect 338172 330500 338580 330528
rect 338172 330488 338178 330500
rect 338574 330488 338580 330500
rect 338632 330488 338638 330540
rect 349982 330488 349988 330540
rect 350040 330528 350046 330540
rect 350442 330528 350448 330540
rect 350040 330500 350448 330528
rect 350040 330488 350046 330500
rect 350442 330488 350448 330500
rect 350500 330488 350506 330540
rect 362402 330488 362408 330540
rect 362460 330528 362466 330540
rect 362862 330528 362868 330540
rect 362460 330500 362868 330528
rect 362460 330488 362466 330500
rect 362862 330488 362868 330500
rect 362920 330488 362926 330540
rect 381354 330488 381360 330540
rect 381412 330528 381418 330540
rect 382090 330528 382096 330540
rect 381412 330500 382096 330528
rect 381412 330488 381418 330500
rect 382090 330488 382096 330500
rect 382148 330488 382154 330540
rect 396350 330488 396356 330540
rect 396408 330528 396414 330540
rect 519538 330528 519544 330540
rect 396408 330500 519544 330528
rect 396408 330488 396414 330500
rect 519538 330488 519544 330500
rect 519596 330488 519602 330540
rect 244458 330460 244464 330472
rect 238726 330432 244464 330460
rect 244458 330420 244464 330432
rect 244516 330420 244522 330472
rect 254026 330420 254032 330472
rect 254084 330460 254090 330472
rect 254946 330460 254952 330472
rect 254084 330432 254952 330460
rect 254084 330420 254090 330432
rect 254946 330420 254952 330432
rect 255004 330420 255010 330472
rect 255406 330420 255412 330472
rect 255464 330460 255470 330472
rect 256050 330460 256056 330472
rect 255464 330432 256056 330460
rect 255464 330420 255470 330432
rect 256050 330420 256056 330432
rect 256108 330420 256114 330472
rect 324406 330420 324412 330472
rect 324464 330460 324470 330472
rect 325418 330460 325424 330472
rect 324464 330432 325424 330460
rect 324464 330420 324470 330432
rect 325418 330420 325424 330432
rect 325476 330420 325482 330472
rect 331306 330420 331312 330472
rect 331364 330460 331370 330472
rect 332318 330460 332324 330472
rect 331364 330432 332324 330460
rect 331364 330420 331370 330432
rect 332318 330420 332324 330432
rect 332376 330420 332382 330472
rect 338206 330420 338212 330472
rect 338264 330460 338270 330472
rect 338942 330460 338948 330472
rect 338264 330432 338948 330460
rect 338264 330420 338270 330432
rect 338942 330420 338948 330432
rect 339000 330420 339006 330472
rect 414290 330420 414296 330472
rect 414348 330460 414354 330472
rect 415118 330460 415124 330472
rect 414348 330432 415124 330460
rect 414348 330420 414354 330432
rect 415118 330420 415124 330432
rect 415176 330420 415182 330472
rect 119982 329332 119988 329384
rect 120040 329372 120046 329384
rect 269114 329372 269120 329384
rect 120040 329344 269120 329372
rect 120040 329332 120046 329344
rect 269114 329332 269120 329344
rect 269172 329332 269178 329384
rect 58618 329264 58624 329316
rect 58676 329304 58682 329316
rect 248690 329304 248696 329316
rect 58676 329276 248696 329304
rect 58676 329264 58682 329276
rect 248690 329264 248696 329276
rect 248748 329264 248754 329316
rect 47578 329196 47584 329248
rect 47636 329236 47642 329248
rect 246574 329236 246580 329248
rect 47636 329208 246580 329236
rect 47636 329196 47642 329208
rect 246574 329196 246580 329208
rect 246632 329196 246638 329248
rect 32398 329128 32404 329180
rect 32456 329168 32462 329180
rect 240318 329168 240324 329180
rect 32456 329140 240324 329168
rect 32456 329128 32462 329140
rect 240318 329128 240324 329140
rect 240376 329128 240382 329180
rect 397362 329128 397368 329180
rect 397420 329168 397426 329180
rect 524414 329168 524420 329180
rect 397420 329140 524420 329168
rect 397420 329128 397426 329140
rect 524414 329128 524420 329140
rect 524472 329128 524478 329180
rect 36538 329060 36544 329112
rect 36596 329100 36602 329112
rect 245654 329100 245660 329112
rect 36596 329072 245660 329100
rect 36596 329060 36602 329072
rect 245654 329060 245660 329072
rect 245712 329060 245718 329112
rect 400766 329060 400772 329112
rect 400824 329100 400830 329112
rect 535454 329100 535460 329112
rect 400824 329072 535460 329100
rect 400824 329060 400830 329072
rect 535454 329060 535460 329072
rect 535512 329060 535518 329112
rect 329834 328040 329840 328092
rect 329892 328080 329898 328092
rect 330570 328080 330576 328092
rect 329892 328052 330576 328080
rect 329892 328040 329898 328052
rect 330570 328040 330576 328052
rect 330628 328040 330634 328092
rect 14458 327700 14464 327752
rect 14516 327740 14522 327752
rect 237742 327740 237748 327752
rect 14516 327712 237748 327740
rect 14516 327700 14522 327712
rect 237742 327700 237748 327712
rect 237800 327700 237806 327752
rect 314746 327156 314752 327208
rect 314804 327196 314810 327208
rect 315574 327196 315580 327208
rect 314804 327168 315580 327196
rect 314804 327156 314810 327168
rect 315574 327156 315580 327168
rect 315632 327156 315638 327208
rect 276198 326408 276204 326460
rect 276256 326408 276262 326460
rect 302510 326448 302516 326460
rect 302471 326420 302516 326448
rect 302510 326408 302516 326420
rect 302568 326408 302574 326460
rect 309226 326408 309232 326460
rect 309284 326448 309290 326460
rect 310054 326448 310060 326460
rect 309284 326420 310060 326448
rect 309284 326408 309290 326420
rect 310054 326408 310060 326420
rect 310112 326408 310118 326460
rect 274726 326340 274732 326392
rect 274784 326380 274790 326392
rect 275738 326380 275744 326392
rect 274784 326352 275744 326380
rect 274784 326340 274790 326352
rect 275738 326340 275744 326352
rect 275796 326340 275802 326392
rect 234706 326272 234712 326324
rect 234764 326312 234770 326324
rect 235534 326312 235540 326324
rect 234764 326284 235540 326312
rect 234764 326272 234770 326284
rect 235534 326272 235540 326284
rect 235592 326272 235598 326324
rect 276216 326256 276244 326408
rect 277486 326340 277492 326392
rect 277544 326380 277550 326392
rect 277670 326380 277676 326392
rect 277544 326352 277676 326380
rect 277544 326340 277550 326352
rect 277670 326340 277676 326352
rect 277728 326340 277734 326392
rect 280246 326340 280252 326392
rect 280304 326380 280310 326392
rect 280890 326380 280896 326392
rect 280304 326352 280896 326380
rect 280304 326340 280310 326352
rect 280890 326340 280896 326352
rect 280948 326340 280954 326392
rect 302326 326340 302332 326392
rect 302384 326380 302390 326392
rect 303154 326380 303160 326392
rect 302384 326352 303160 326380
rect 302384 326340 302390 326352
rect 303154 326340 303160 326352
rect 303212 326340 303218 326392
rect 304994 326340 305000 326392
rect 305052 326380 305058 326392
rect 305362 326380 305368 326392
rect 305052 326352 305368 326380
rect 305052 326340 305058 326352
rect 305362 326340 305368 326352
rect 305420 326340 305426 326392
rect 306374 326340 306380 326392
rect 306432 326380 306438 326392
rect 307478 326380 307484 326392
rect 306432 326352 307484 326380
rect 306432 326340 306438 326352
rect 307478 326340 307484 326352
rect 307536 326340 307542 326392
rect 307754 326340 307760 326392
rect 307812 326380 307818 326392
rect 308582 326380 308588 326392
rect 307812 326352 308588 326380
rect 307812 326340 307818 326352
rect 308582 326340 308588 326352
rect 308640 326340 308646 326392
rect 309134 326340 309140 326392
rect 309192 326380 309198 326392
rect 309686 326380 309692 326392
rect 309192 326352 309692 326380
rect 309192 326340 309198 326352
rect 309686 326340 309692 326352
rect 309744 326340 309750 326392
rect 310606 326340 310612 326392
rect 310664 326380 310670 326392
rect 311158 326380 311164 326392
rect 310664 326352 311164 326380
rect 310664 326340 310670 326352
rect 311158 326340 311164 326352
rect 311216 326340 311222 326392
rect 276198 326204 276204 326256
rect 276256 326204 276262 326256
rect 277486 326204 277492 326256
rect 277544 326244 277550 326256
rect 278314 326244 278320 326256
rect 277544 326216 278320 326244
rect 277544 326204 277550 326216
rect 278314 326204 278320 326216
rect 278372 326204 278378 326256
rect 305086 326204 305092 326256
rect 305144 326244 305150 326256
rect 305730 326244 305736 326256
rect 305144 326216 305736 326244
rect 305144 326204 305150 326216
rect 305730 326204 305736 326216
rect 305788 326204 305794 326256
rect 305178 326136 305184 326188
rect 305236 326176 305242 326188
rect 306098 326176 306104 326188
rect 305236 326148 306104 326176
rect 305236 326136 305242 326148
rect 306098 326136 306104 326148
rect 306156 326136 306162 326188
rect 421650 325592 421656 325644
rect 421708 325632 421714 325644
rect 579890 325632 579896 325644
rect 421708 325604 579896 325632
rect 421708 325592 421714 325604
rect 579890 325592 579896 325604
rect 579948 325592 579954 325644
rect 302510 323592 302516 323604
rect 302471 323564 302516 323592
rect 302510 323552 302516 323564
rect 302568 323552 302574 323604
rect 276106 321512 276112 321564
rect 276164 321552 276170 321564
rect 276290 321552 276296 321564
rect 276164 321524 276296 321552
rect 276164 321512 276170 321524
rect 276290 321512 276296 321524
rect 276348 321512 276354 321564
rect 555418 313216 555424 313268
rect 555476 313256 555482 313268
rect 580166 313256 580172 313268
rect 555476 313228 580172 313256
rect 555476 313216 555482 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 232590 215268 232596 215280
rect 3384 215240 232596 215268
rect 3384 215228 3390 215240
rect 232590 215228 232596 215240
rect 232648 215228 232654 215280
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 226978 45540 226984 45552
rect 3476 45512 226984 45540
rect 3476 45500 3482 45512
rect 226978 45500 226984 45512
rect 227036 45500 227042 45552
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 414934 20652 414940 20664
rect 3476 20624 414940 20652
rect 3476 20612 3482 20624
rect 414934 20612 414940 20624
rect 414992 20612 414998 20664
rect 431218 20612 431224 20664
rect 431276 20652 431282 20664
rect 579982 20652 579988 20664
rect 431276 20624 579988 20652
rect 431276 20612 431282 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 157242 18572 157248 18624
rect 157300 18612 157306 18624
rect 282178 18612 282184 18624
rect 157300 18584 282184 18612
rect 157300 18572 157306 18584
rect 282178 18572 282184 18584
rect 282236 18572 282242 18624
rect 161290 17212 161296 17264
rect 161348 17252 161354 17264
rect 284386 17252 284392 17264
rect 161348 17224 284392 17252
rect 161348 17212 161354 17224
rect 284386 17212 284392 17224
rect 284444 17212 284450 17264
rect 139302 15852 139308 15904
rect 139360 15892 139366 15904
rect 277578 15892 277584 15904
rect 139360 15864 277584 15892
rect 139360 15852 139366 15864
rect 277578 15852 277584 15864
rect 277636 15852 277642 15904
rect 252370 14424 252376 14476
rect 252428 14464 252434 14476
rect 311986 14464 311992 14476
rect 252428 14436 311992 14464
rect 252428 14424 252434 14436
rect 311986 14424 311992 14436
rect 312044 14424 312050 14476
rect 184934 13336 184940 13388
rect 184992 13376 184998 13388
rect 291286 13376 291292 13388
rect 184992 13348 291292 13376
rect 184992 13336 184998 13348
rect 291286 13336 291292 13348
rect 291344 13336 291350 13388
rect 125870 13268 125876 13320
rect 125928 13308 125934 13320
rect 233970 13308 233976 13320
rect 125928 13280 233976 13308
rect 125928 13268 125934 13280
rect 233970 13268 233976 13280
rect 234028 13268 234034 13320
rect 164142 13200 164148 13252
rect 164200 13240 164206 13252
rect 284478 13240 284484 13252
rect 164200 13212 284484 13240
rect 164200 13200 164206 13212
rect 284478 13200 284484 13212
rect 284536 13200 284542 13252
rect 149974 13132 149980 13184
rect 150032 13172 150038 13184
rect 280246 13172 280252 13184
rect 150032 13144 280252 13172
rect 150032 13132 150038 13144
rect 280246 13132 280252 13144
rect 280304 13132 280310 13184
rect 128170 13064 128176 13116
rect 128228 13104 128234 13116
rect 273438 13104 273444 13116
rect 128228 13076 273444 13104
rect 128228 13064 128234 13076
rect 273438 13064 273444 13076
rect 273496 13064 273502 13116
rect 212166 12180 212172 12232
rect 212224 12220 212230 12232
rect 233878 12220 233884 12232
rect 212224 12192 233884 12220
rect 212224 12180 212230 12192
rect 233878 12180 233884 12192
rect 233936 12180 233942 12232
rect 182542 12112 182548 12164
rect 182600 12152 182606 12164
rect 224218 12152 224224 12164
rect 182600 12124 224224 12152
rect 182600 12112 182606 12124
rect 224218 12112 224224 12124
rect 224276 12112 224282 12164
rect 175918 12044 175924 12096
rect 175976 12084 175982 12096
rect 228358 12084 228364 12096
rect 175976 12056 228364 12084
rect 175976 12044 175982 12056
rect 228358 12044 228364 12056
rect 228416 12044 228422 12096
rect 164878 11976 164884 12028
rect 164936 12016 164942 12028
rect 231118 12016 231124 12028
rect 164936 11988 231124 12016
rect 164936 11976 164942 11988
rect 231118 11976 231124 11988
rect 231176 11976 231182 12028
rect 154206 11908 154212 11960
rect 154264 11948 154270 11960
rect 232498 11948 232504 11960
rect 154264 11920 232504 11948
rect 154264 11908 154270 11920
rect 232498 11908 232504 11920
rect 232556 11908 232562 11960
rect 251082 11908 251088 11960
rect 251140 11948 251146 11960
rect 291838 11948 291844 11960
rect 251140 11920 291844 11948
rect 251140 11908 251146 11920
rect 291838 11908 291844 11920
rect 291896 11908 291902 11960
rect 167638 11840 167644 11892
rect 167696 11880 167702 11892
rect 285766 11880 285772 11892
rect 167696 11852 285772 11880
rect 167696 11840 167702 11852
rect 285766 11840 285772 11852
rect 285824 11840 285830 11892
rect 78582 11772 78588 11824
rect 78640 11812 78646 11824
rect 258350 11812 258356 11824
rect 78640 11784 258356 11812
rect 78640 11772 78646 11784
rect 258350 11772 258356 11784
rect 258408 11772 258414 11824
rect 74442 11704 74448 11756
rect 74500 11744 74506 11756
rect 256878 11744 256884 11756
rect 74500 11716 256884 11744
rect 74500 11704 74506 11716
rect 256878 11704 256884 11716
rect 256936 11704 256942 11756
rect 440326 11704 440332 11756
rect 440384 11744 440390 11756
rect 441522 11744 441528 11756
rect 440384 11716 441528 11744
rect 440384 11704 440390 11716
rect 441522 11704 441528 11716
rect 441580 11704 441586 11756
rect 448606 11704 448612 11756
rect 448664 11744 448670 11756
rect 449802 11744 449808 11756
rect 448664 11716 449808 11744
rect 448664 11704 448670 11716
rect 449802 11704 449808 11716
rect 449860 11704 449866 11756
rect 160094 11636 160100 11688
rect 160152 11676 160158 11688
rect 161290 11676 161296 11688
rect 160152 11648 161296 11676
rect 160152 11636 160158 11648
rect 161290 11636 161296 11648
rect 161348 11636 161354 11688
rect 95050 10956 95056 11008
rect 95108 10996 95114 11008
rect 263686 10996 263692 11008
rect 95108 10968 263692 10996
rect 95108 10956 95114 10968
rect 263686 10956 263692 10968
rect 263744 10956 263750 11008
rect 428458 10956 428464 11008
rect 428516 10996 428522 11008
rect 430850 10996 430856 11008
rect 428516 10968 430856 10996
rect 428516 10956 428522 10968
rect 430850 10956 430856 10968
rect 430908 10956 430914 11008
rect 91002 10888 91008 10940
rect 91060 10928 91066 10940
rect 262398 10928 262404 10940
rect 91060 10900 262404 10928
rect 91060 10888 91066 10900
rect 262398 10888 262404 10900
rect 262456 10888 262462 10940
rect 70302 10820 70308 10872
rect 70360 10860 70366 10872
rect 255590 10860 255596 10872
rect 70360 10832 255596 10860
rect 70360 10820 70366 10832
rect 255590 10820 255596 10832
rect 255648 10820 255654 10872
rect 67542 10752 67548 10804
rect 67600 10792 67606 10804
rect 255498 10792 255504 10804
rect 67600 10764 255504 10792
rect 67600 10752 67606 10764
rect 255498 10752 255504 10764
rect 255556 10752 255562 10804
rect 63218 10684 63224 10736
rect 63276 10724 63282 10736
rect 254210 10724 254216 10736
rect 63276 10696 254216 10724
rect 63276 10684 63282 10696
rect 254210 10684 254216 10696
rect 254268 10684 254274 10736
rect 60642 10616 60648 10668
rect 60700 10656 60706 10668
rect 252738 10656 252744 10668
rect 60700 10628 252744 10656
rect 60700 10616 60706 10628
rect 252738 10616 252744 10628
rect 252796 10616 252802 10668
rect 260650 10616 260656 10668
rect 260708 10656 260714 10668
rect 286318 10656 286324 10668
rect 260708 10628 286324 10656
rect 260708 10616 260714 10628
rect 286318 10616 286324 10628
rect 286376 10616 286382 10668
rect 56502 10548 56508 10600
rect 56560 10588 56566 10600
rect 251266 10588 251272 10600
rect 56560 10560 251272 10588
rect 56560 10548 56566 10560
rect 251266 10548 251272 10560
rect 251324 10548 251330 10600
rect 253842 10548 253848 10600
rect 253900 10588 253906 10600
rect 289078 10588 289084 10600
rect 253900 10560 289084 10588
rect 253900 10548 253906 10560
rect 289078 10548 289084 10560
rect 289136 10548 289142 10600
rect 53742 10480 53748 10532
rect 53800 10520 53806 10532
rect 249978 10520 249984 10532
rect 53800 10492 249984 10520
rect 53800 10480 53806 10492
rect 249978 10480 249984 10492
rect 250036 10480 250042 10532
rect 271782 10480 271788 10532
rect 271840 10520 271846 10532
rect 317598 10520 317604 10532
rect 271840 10492 317604 10520
rect 271840 10480 271846 10492
rect 317598 10480 317604 10492
rect 317656 10480 317662 10532
rect 49602 10412 49608 10464
rect 49660 10452 49666 10464
rect 249886 10452 249892 10464
rect 49660 10424 249892 10452
rect 49660 10412 49666 10424
rect 249886 10412 249892 10424
rect 249944 10412 249950 10464
rect 269022 10412 269028 10464
rect 269080 10452 269086 10464
rect 317506 10452 317512 10464
rect 269080 10424 317512 10452
rect 269080 10412 269086 10424
rect 317506 10412 317512 10424
rect 317564 10412 317570 10464
rect 45462 10344 45468 10396
rect 45520 10384 45526 10396
rect 248598 10384 248604 10396
rect 45520 10356 248604 10384
rect 45520 10344 45526 10356
rect 248598 10344 248604 10356
rect 248656 10344 248662 10396
rect 264882 10344 264888 10396
rect 264940 10384 264946 10396
rect 316126 10384 316132 10396
rect 264940 10356 316132 10384
rect 264940 10344 264946 10356
rect 316126 10344 316132 10356
rect 316184 10344 316190 10396
rect 41322 10276 41328 10328
rect 41380 10316 41386 10328
rect 247126 10316 247132 10328
rect 41380 10288 247132 10316
rect 41380 10276 41386 10288
rect 247126 10276 247132 10288
rect 247184 10276 247190 10328
rect 256602 10276 256608 10328
rect 256660 10316 256666 10328
rect 313458 10316 313464 10328
rect 256660 10288 313464 10316
rect 256660 10276 256666 10288
rect 313458 10276 313464 10288
rect 313516 10276 313522 10328
rect 357158 10276 357164 10328
rect 357216 10316 357222 10328
rect 392578 10316 392584 10328
rect 357216 10288 392584 10316
rect 357216 10276 357222 10288
rect 392578 10276 392584 10288
rect 392636 10276 392642 10328
rect 97902 10208 97908 10260
rect 97960 10248 97966 10260
rect 265066 10248 265072 10260
rect 97960 10220 265072 10248
rect 97960 10208 97966 10220
rect 265066 10208 265072 10220
rect 265124 10208 265130 10260
rect 102042 10140 102048 10192
rect 102100 10180 102106 10192
rect 265158 10180 265164 10192
rect 102100 10152 265164 10180
rect 102100 10140 102106 10152
rect 265158 10140 265164 10152
rect 265216 10140 265222 10192
rect 104526 10072 104532 10124
rect 104584 10112 104590 10124
rect 266446 10112 266452 10124
rect 104584 10084 266452 10112
rect 104584 10072 104590 10084
rect 266446 10072 266452 10084
rect 266504 10072 266510 10124
rect 108942 10004 108948 10056
rect 109000 10044 109006 10056
rect 267826 10044 267832 10056
rect 109000 10016 267832 10044
rect 109000 10004 109006 10016
rect 267826 10004 267832 10016
rect 267884 10004 267890 10056
rect 111610 9936 111616 9988
rect 111668 9976 111674 9988
rect 269298 9976 269304 9988
rect 111668 9948 269304 9976
rect 111668 9936 111674 9948
rect 269298 9936 269304 9948
rect 269356 9936 269362 9988
rect 115842 9868 115848 9920
rect 115900 9908 115906 9920
rect 270678 9908 270684 9920
rect 115900 9880 270684 9908
rect 115900 9868 115906 9880
rect 270678 9868 270684 9880
rect 270736 9868 270742 9920
rect 119798 9800 119804 9852
rect 119856 9840 119862 9852
rect 270586 9840 270592 9852
rect 119856 9812 270592 9840
rect 119856 9800 119862 9812
rect 270586 9800 270592 9812
rect 270644 9800 270650 9852
rect 122742 9732 122748 9784
rect 122800 9772 122806 9784
rect 271966 9772 271972 9784
rect 122800 9744 271972 9772
rect 122800 9732 122806 9744
rect 271966 9732 271972 9744
rect 272024 9732 272030 9784
rect 209774 9596 209780 9648
rect 209832 9636 209838 9648
rect 299658 9636 299664 9648
rect 209832 9608 299664 9636
rect 209832 9596 209838 9608
rect 299658 9596 299664 9608
rect 299716 9596 299722 9648
rect 417510 9596 417516 9648
rect 417568 9636 417574 9648
rect 420178 9636 420184 9648
rect 417568 9608 420184 9636
rect 417568 9596 417574 9608
rect 420178 9596 420184 9608
rect 420236 9596 420242 9648
rect 206186 9528 206192 9580
rect 206244 9568 206250 9580
rect 298186 9568 298192 9580
rect 206244 9540 298192 9568
rect 206244 9528 206250 9540
rect 298186 9528 298192 9540
rect 298244 9528 298250 9580
rect 202690 9460 202696 9512
rect 202748 9500 202754 9512
rect 296806 9500 296812 9512
rect 202748 9472 296812 9500
rect 202748 9460 202754 9472
rect 296806 9460 296812 9472
rect 296864 9460 296870 9512
rect 199102 9392 199108 9444
rect 199160 9432 199166 9444
rect 295518 9432 295524 9444
rect 199160 9404 295524 9432
rect 199160 9392 199166 9404
rect 295518 9392 295524 9404
rect 295576 9392 295582 9444
rect 195606 9324 195612 9376
rect 195664 9364 195670 9376
rect 294138 9364 294144 9376
rect 195664 9336 294144 9364
rect 195664 9324 195670 9336
rect 294138 9324 294144 9336
rect 294196 9324 294202 9376
rect 192018 9256 192024 9308
rect 192076 9296 192082 9308
rect 294046 9296 294052 9308
rect 192076 9268 294052 9296
rect 192076 9256 192082 9268
rect 294046 9256 294052 9268
rect 294104 9256 294110 9308
rect 135254 9188 135260 9240
rect 135312 9228 135318 9240
rect 276106 9228 276112 9240
rect 135312 9200 276112 9228
rect 135312 9188 135318 9200
rect 276106 9188 276112 9200
rect 276164 9188 276170 9240
rect 131758 9120 131764 9172
rect 131816 9160 131822 9172
rect 274910 9160 274916 9172
rect 131816 9132 274916 9160
rect 131816 9120 131822 9132
rect 274910 9120 274916 9132
rect 274968 9120 274974 9172
rect 37182 9052 37188 9104
rect 37240 9092 37246 9104
rect 245930 9092 245936 9104
rect 37240 9064 245936 9092
rect 37240 9052 37246 9064
rect 245930 9052 245936 9064
rect 245988 9052 245994 9104
rect 248782 9052 248788 9104
rect 248840 9092 248846 9104
rect 310790 9092 310796 9104
rect 248840 9064 310796 9092
rect 248840 9052 248846 9064
rect 310790 9052 310796 9064
rect 310848 9052 310854 9104
rect 418798 9052 418804 9104
rect 418856 9092 418862 9104
rect 427262 9092 427268 9104
rect 418856 9064 427268 9092
rect 418856 9052 418862 9064
rect 427262 9052 427268 9064
rect 427320 9052 427326 9104
rect 33594 8984 33600 9036
rect 33652 9024 33658 9036
rect 244366 9024 244372 9036
rect 33652 8996 244372 9024
rect 33652 8984 33658 8996
rect 244366 8984 244372 8996
rect 244424 8984 244430 9036
rect 245194 8984 245200 9036
rect 245252 9024 245258 9036
rect 310698 9024 310704 9036
rect 245252 8996 310704 9024
rect 245252 8984 245258 8996
rect 310698 8984 310704 8996
rect 310756 8984 310762 9036
rect 353938 8984 353944 9036
rect 353996 9024 354002 9036
rect 370590 9024 370596 9036
rect 353996 8996 370596 9024
rect 353996 8984 354002 8996
rect 370590 8984 370596 8996
rect 370648 8984 370654 9036
rect 372430 8984 372436 9036
rect 372488 9024 372494 9036
rect 445018 9024 445024 9036
rect 372488 8996 445024 9024
rect 372488 8984 372494 8996
rect 445018 8984 445024 8996
rect 445076 8984 445082 9036
rect 8754 8916 8760 8968
rect 8812 8956 8818 8968
rect 237466 8956 237472 8968
rect 8812 8928 237472 8956
rect 8812 8916 8818 8928
rect 237466 8916 237472 8928
rect 237524 8916 237530 8968
rect 238110 8916 238116 8968
rect 238168 8956 238174 8968
rect 307938 8956 307944 8968
rect 238168 8928 307944 8956
rect 238168 8916 238174 8928
rect 307938 8916 307944 8928
rect 307996 8916 308002 8968
rect 353018 8916 353024 8968
rect 353076 8956 353082 8968
rect 382366 8956 382372 8968
rect 353076 8928 382372 8956
rect 353076 8916 353082 8928
rect 382366 8916 382372 8928
rect 382424 8916 382430 8968
rect 382918 8916 382924 8968
rect 382976 8956 382982 8968
rect 416682 8956 416688 8968
rect 382976 8928 416688 8956
rect 382976 8916 382982 8928
rect 416682 8916 416688 8928
rect 416740 8916 416746 8968
rect 417418 8916 417424 8968
rect 417476 8956 417482 8968
rect 494698 8956 494704 8968
rect 417476 8928 494704 8956
rect 417476 8916 417482 8928
rect 494698 8916 494704 8928
rect 494756 8916 494762 8968
rect 126974 8848 126980 8900
rect 127032 8888 127038 8900
rect 213178 8888 213184 8900
rect 127032 8860 213184 8888
rect 127032 8848 127038 8860
rect 213178 8848 213184 8860
rect 213236 8848 213242 8900
rect 213362 8848 213368 8900
rect 213420 8888 213426 8900
rect 299566 8888 299572 8900
rect 213420 8860 299572 8888
rect 213420 8848 213426 8860
rect 299566 8848 299572 8860
rect 299624 8848 299630 8900
rect 216858 8780 216864 8832
rect 216916 8820 216922 8832
rect 300946 8820 300952 8832
rect 216916 8792 300952 8820
rect 216916 8780 216922 8792
rect 300946 8780 300952 8792
rect 301004 8780 301010 8832
rect 220446 8712 220452 8764
rect 220504 8752 220510 8764
rect 302418 8752 302424 8764
rect 220504 8724 302424 8752
rect 220504 8712 220510 8724
rect 302418 8712 302424 8724
rect 302476 8712 302482 8764
rect 223942 8644 223948 8696
rect 224000 8684 224006 8696
rect 303706 8684 303712 8696
rect 224000 8656 303712 8684
rect 224000 8644 224006 8656
rect 303706 8644 303712 8656
rect 303764 8644 303770 8696
rect 227530 8576 227536 8628
rect 227588 8616 227594 8628
rect 305270 8616 305276 8628
rect 227588 8588 305276 8616
rect 227588 8576 227594 8588
rect 305270 8576 305276 8588
rect 305328 8576 305334 8628
rect 231026 8508 231032 8560
rect 231084 8548 231090 8560
rect 305178 8548 305184 8560
rect 231084 8520 305184 8548
rect 231084 8508 231090 8520
rect 305178 8508 305184 8520
rect 305236 8508 305242 8560
rect 234982 8440 234988 8492
rect 235040 8480 235046 8492
rect 306650 8480 306656 8492
rect 235040 8452 306656 8480
rect 235040 8440 235046 8452
rect 306650 8440 306656 8452
rect 306708 8440 306714 8492
rect 241698 8372 241704 8424
rect 241756 8412 241762 8424
rect 309410 8412 309416 8424
rect 241756 8384 309416 8412
rect 241756 8372 241762 8384
rect 309410 8372 309416 8384
rect 309468 8372 309474 8424
rect 421558 8304 421564 8356
rect 421616 8344 421622 8356
rect 423766 8344 423772 8356
rect 421616 8316 423772 8344
rect 421616 8304 421622 8316
rect 423766 8304 423772 8316
rect 423824 8304 423830 8356
rect 137646 8236 137652 8288
rect 137704 8276 137710 8288
rect 277670 8276 277676 8288
rect 137704 8248 277676 8276
rect 137704 8236 137710 8248
rect 277670 8236 277676 8248
rect 277728 8236 277734 8288
rect 372338 8236 372344 8288
rect 372396 8276 372402 8288
rect 442626 8276 442632 8288
rect 372396 8248 442632 8276
rect 372396 8236 372402 8248
rect 442626 8236 442632 8248
rect 442684 8236 442690 8288
rect 134150 8168 134156 8220
rect 134208 8208 134214 8220
rect 276198 8208 276204 8220
rect 134208 8180 276204 8208
rect 134208 8168 134214 8180
rect 276198 8168 276204 8180
rect 276256 8168 276262 8220
rect 403986 8168 403992 8220
rect 404044 8208 404050 8220
rect 545482 8208 545488 8220
rect 404044 8180 545488 8208
rect 404044 8168 404050 8180
rect 545482 8168 545488 8180
rect 545540 8168 545546 8220
rect 79686 8100 79692 8152
rect 79744 8140 79750 8152
rect 258077 8143 258135 8149
rect 258077 8140 258089 8143
rect 79744 8112 258089 8140
rect 79744 8100 79750 8112
rect 258077 8109 258089 8112
rect 258123 8109 258135 8143
rect 258350 8140 258356 8152
rect 258077 8103 258135 8109
rect 258184 8112 258356 8140
rect 76190 8032 76196 8084
rect 76248 8072 76254 8084
rect 258184 8072 258212 8112
rect 258350 8100 258356 8112
rect 258408 8100 258414 8152
rect 258445 8143 258503 8149
rect 258445 8109 258457 8143
rect 258491 8140 258503 8143
rect 259546 8140 259552 8152
rect 258491 8112 259552 8140
rect 258491 8109 258503 8112
rect 258445 8103 258503 8109
rect 259546 8100 259552 8112
rect 259604 8100 259610 8152
rect 265342 8100 265348 8152
rect 265400 8140 265406 8152
rect 316218 8140 316224 8152
rect 265400 8112 316224 8140
rect 265400 8100 265406 8112
rect 316218 8100 316224 8112
rect 316276 8100 316282 8152
rect 405366 8100 405372 8152
rect 405424 8140 405430 8152
rect 549070 8140 549076 8152
rect 405424 8112 549076 8140
rect 405424 8100 405430 8112
rect 549070 8100 549076 8112
rect 549128 8100 549134 8152
rect 76248 8044 258212 8072
rect 76248 8032 76254 8044
rect 258258 8032 258264 8084
rect 258316 8072 258322 8084
rect 258316 8044 261064 8072
rect 258316 8032 258322 8044
rect 72602 7964 72608 8016
rect 72660 8004 72666 8016
rect 256786 8004 256792 8016
rect 72660 7976 256792 8004
rect 72660 7964 72666 7976
rect 256786 7964 256792 7976
rect 256844 7964 256850 8016
rect 258077 8007 258135 8013
rect 258077 7973 258089 8007
rect 258123 8004 258135 8007
rect 261036 8004 261064 8044
rect 261754 8032 261760 8084
rect 261812 8072 261818 8084
rect 314746 8072 314752 8084
rect 261812 8044 314752 8072
rect 261812 8032 261818 8044
rect 314746 8032 314752 8044
rect 314804 8032 314810 8084
rect 405458 8032 405464 8084
rect 405516 8072 405522 8084
rect 552658 8072 552664 8084
rect 405516 8044 552664 8072
rect 405516 8032 405522 8044
rect 552658 8032 552664 8044
rect 552716 8032 552722 8084
rect 314838 8004 314844 8016
rect 258123 7976 258304 8004
rect 261036 7976 314844 8004
rect 258123 7973 258135 7976
rect 258077 7967 258135 7973
rect 30098 7896 30104 7948
rect 30156 7936 30162 7948
rect 243078 7936 243084 7948
rect 30156 7908 243084 7936
rect 30156 7896 30162 7908
rect 243078 7896 243084 7908
rect 243136 7896 243142 7948
rect 251174 7896 251180 7948
rect 251232 7936 251238 7948
rect 258276 7936 258304 7976
rect 314838 7964 314844 7976
rect 314896 7964 314902 8016
rect 406746 7964 406752 8016
rect 406804 8004 406810 8016
rect 556154 8004 556160 8016
rect 406804 7976 556160 8004
rect 406804 7964 406810 7976
rect 556154 7964 556160 7976
rect 556212 7964 556218 8016
rect 313366 7936 313372 7948
rect 251232 7908 258212 7936
rect 258276 7908 313372 7936
rect 251232 7896 251238 7908
rect 26510 7828 26516 7880
rect 26568 7868 26574 7880
rect 242986 7868 242992 7880
rect 26568 7840 242992 7868
rect 26568 7828 26574 7840
rect 242986 7828 242992 7840
rect 243044 7828 243050 7880
rect 254670 7828 254676 7880
rect 254728 7868 254734 7880
rect 258077 7871 258135 7877
rect 258077 7868 258089 7871
rect 254728 7840 258089 7868
rect 254728 7828 254734 7840
rect 258077 7837 258089 7840
rect 258123 7837 258135 7871
rect 258184 7868 258212 7908
rect 313366 7896 313372 7908
rect 313424 7896 313430 7948
rect 408218 7896 408224 7948
rect 408276 7936 408282 7948
rect 559742 7936 559748 7948
rect 408276 7908 559748 7936
rect 408276 7896 408282 7908
rect 559742 7896 559748 7908
rect 559800 7896 559806 7948
rect 312078 7868 312084 7880
rect 258184 7840 312084 7868
rect 258077 7831 258135 7837
rect 312078 7828 312084 7840
rect 312136 7828 312142 7880
rect 409506 7828 409512 7880
rect 409564 7868 409570 7880
rect 563238 7868 563244 7880
rect 409564 7840 563244 7868
rect 409564 7828 409570 7840
rect 563238 7828 563244 7840
rect 563296 7828 563302 7880
rect 21818 7760 21824 7812
rect 21876 7800 21882 7812
rect 241790 7800 241796 7812
rect 21876 7772 241796 7800
rect 21876 7760 21882 7772
rect 241790 7760 241796 7772
rect 241848 7760 241854 7812
rect 247586 7760 247592 7812
rect 247644 7800 247650 7812
rect 310606 7800 310612 7812
rect 247644 7772 310612 7800
rect 247644 7760 247650 7772
rect 310606 7760 310612 7772
rect 310664 7760 310670 7812
rect 410978 7760 410984 7812
rect 411036 7800 411042 7812
rect 566826 7800 566832 7812
rect 411036 7772 566832 7800
rect 411036 7760 411042 7772
rect 566826 7760 566832 7772
rect 566884 7760 566890 7812
rect 17034 7692 17040 7744
rect 17092 7732 17098 7744
rect 240134 7732 240140 7744
rect 17092 7704 240140 7732
rect 17092 7692 17098 7704
rect 240134 7692 240140 7704
rect 240192 7692 240198 7744
rect 244090 7692 244096 7744
rect 244148 7732 244154 7744
rect 309226 7732 309232 7744
rect 244148 7704 309232 7732
rect 244148 7692 244154 7704
rect 309226 7692 309232 7704
rect 309284 7692 309290 7744
rect 410886 7692 410892 7744
rect 410944 7732 410950 7744
rect 570322 7732 570328 7744
rect 410944 7704 570328 7732
rect 410944 7692 410950 7704
rect 570322 7692 570328 7704
rect 570380 7692 570386 7744
rect 12342 7624 12348 7676
rect 12400 7664 12406 7676
rect 237374 7664 237380 7676
rect 12400 7636 237380 7664
rect 12400 7624 12406 7636
rect 237374 7624 237380 7636
rect 237432 7624 237438 7676
rect 240502 7624 240508 7676
rect 240560 7664 240566 7676
rect 309318 7664 309324 7676
rect 240560 7636 309324 7664
rect 240560 7624 240566 7636
rect 309318 7624 309324 7636
rect 309376 7624 309382 7676
rect 412266 7624 412272 7676
rect 412324 7664 412330 7676
rect 573910 7664 573916 7676
rect 412324 7636 573916 7664
rect 412324 7624 412330 7636
rect 573910 7624 573916 7636
rect 573968 7624 573974 7676
rect 4062 7556 4068 7608
rect 4120 7596 4126 7608
rect 236178 7596 236184 7608
rect 4120 7568 236184 7596
rect 4120 7556 4126 7568
rect 236178 7556 236184 7568
rect 236236 7556 236242 7608
rect 237006 7556 237012 7608
rect 237064 7596 237070 7608
rect 307846 7596 307852 7608
rect 237064 7568 307852 7596
rect 237064 7556 237070 7568
rect 307846 7556 307852 7568
rect 307904 7556 307910 7608
rect 413738 7556 413744 7608
rect 413796 7596 413802 7608
rect 577406 7596 577412 7608
rect 413796 7568 577412 7596
rect 413796 7556 413802 7568
rect 577406 7556 577412 7568
rect 577464 7556 577470 7608
rect 141234 7488 141240 7540
rect 141292 7528 141298 7540
rect 277486 7528 277492 7540
rect 141292 7500 277492 7528
rect 141292 7488 141298 7500
rect 277486 7488 277492 7500
rect 277544 7488 277550 7540
rect 371050 7488 371056 7540
rect 371108 7528 371114 7540
rect 371108 7500 432552 7528
rect 371108 7488 371114 7500
rect 144730 7420 144736 7472
rect 144788 7460 144794 7472
rect 278958 7460 278964 7472
rect 144788 7432 278964 7460
rect 144788 7420 144794 7432
rect 278958 7420 278964 7432
rect 279016 7420 279022 7472
rect 369670 7420 369676 7472
rect 369728 7460 369734 7472
rect 369728 7432 432460 7460
rect 369728 7420 369734 7432
rect 148318 7352 148324 7404
rect 148376 7392 148382 7404
rect 280338 7392 280344 7404
rect 148376 7364 280344 7392
rect 148376 7352 148382 7364
rect 280338 7352 280344 7364
rect 280396 7352 280402 7404
rect 368382 7352 368388 7404
rect 368440 7392 368446 7404
rect 432046 7392 432052 7404
rect 368440 7364 432052 7392
rect 368440 7352 368446 7364
rect 432046 7352 432052 7364
rect 432104 7352 432110 7404
rect 151814 7284 151820 7336
rect 151872 7324 151878 7336
rect 281718 7324 281724 7336
rect 151872 7296 281724 7324
rect 151872 7284 151878 7296
rect 281718 7284 281724 7296
rect 281776 7284 281782 7336
rect 368290 7284 368296 7336
rect 368348 7324 368354 7336
rect 428458 7324 428464 7336
rect 368348 7296 428464 7324
rect 368348 7284 368354 7296
rect 428458 7284 428464 7296
rect 428516 7284 428522 7336
rect 432432 7324 432460 7432
rect 432524 7392 432552 7500
rect 432598 7488 432604 7540
rect 432656 7528 432662 7540
rect 434438 7528 434444 7540
rect 432656 7500 434444 7528
rect 432656 7488 432662 7500
rect 434438 7488 434444 7500
rect 434496 7488 434502 7540
rect 435358 7488 435364 7540
rect 435416 7528 435422 7540
rect 437934 7528 437940 7540
rect 435416 7500 437940 7528
rect 435416 7488 435422 7500
rect 437934 7488 437940 7500
rect 437992 7488 437998 7540
rect 439130 7392 439136 7404
rect 432524 7364 439136 7392
rect 439130 7352 439136 7364
rect 439188 7352 439194 7404
rect 435542 7324 435548 7336
rect 432432 7296 435548 7324
rect 435542 7284 435548 7296
rect 435600 7284 435606 7336
rect 155402 7216 155408 7268
rect 155460 7256 155466 7268
rect 283006 7256 283012 7268
rect 155460 7228 283012 7256
rect 155460 7216 155466 7228
rect 283006 7216 283012 7228
rect 283064 7216 283070 7268
rect 367002 7216 367008 7268
rect 367060 7256 367066 7268
rect 424962 7256 424968 7268
rect 367060 7228 424968 7256
rect 367060 7216 367066 7228
rect 424962 7216 424968 7228
rect 425020 7216 425026 7268
rect 158898 7148 158904 7200
rect 158956 7188 158962 7200
rect 283098 7188 283104 7200
rect 158956 7160 283104 7188
rect 158956 7148 158962 7160
rect 283098 7148 283104 7160
rect 283156 7148 283162 7200
rect 365530 7148 365536 7200
rect 365588 7188 365594 7200
rect 421374 7188 421380 7200
rect 365588 7160 421380 7188
rect 365588 7148 365594 7160
rect 421374 7148 421380 7160
rect 421432 7148 421438 7200
rect 229830 7080 229836 7132
rect 229888 7120 229894 7132
rect 305086 7120 305092 7132
rect 229888 7092 305092 7120
rect 229888 7080 229894 7092
rect 305086 7080 305092 7092
rect 305144 7080 305150 7132
rect 364150 7080 364156 7132
rect 364208 7120 364214 7132
rect 417878 7120 417884 7132
rect 364208 7092 417884 7120
rect 364208 7080 364214 7092
rect 417878 7080 417884 7092
rect 417936 7080 417942 7132
rect 233418 7012 233424 7064
rect 233476 7052 233482 7064
rect 306558 7052 306564 7064
rect 233476 7024 306564 7052
rect 233476 7012 233482 7024
rect 306558 7012 306564 7024
rect 306616 7012 306622 7064
rect 362586 7012 362592 7064
rect 362644 7052 362650 7064
rect 414290 7052 414296 7064
rect 362644 7024 414296 7052
rect 362644 7012 362650 7024
rect 414290 7012 414296 7024
rect 414348 7012 414354 7064
rect 234614 6808 234620 6860
rect 234672 6848 234678 6860
rect 580166 6848 580172 6860
rect 234672 6820 580172 6848
rect 234672 6808 234678 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 169570 6740 169576 6792
rect 169628 6780 169634 6792
rect 287238 6780 287244 6792
rect 169628 6752 287244 6780
rect 169628 6740 169634 6752
rect 287238 6740 287244 6752
rect 287296 6740 287302 6792
rect 381998 6740 382004 6792
rect 382056 6780 382062 6792
rect 476942 6780 476948 6792
rect 382056 6752 476948 6780
rect 382056 6740 382062 6752
rect 476942 6740 476948 6752
rect 477000 6740 477006 6792
rect 166074 6672 166080 6724
rect 166132 6712 166138 6724
rect 285858 6712 285864 6724
rect 166132 6684 285864 6712
rect 166132 6672 166138 6684
rect 285858 6672 285864 6684
rect 285916 6672 285922 6724
rect 384850 6672 384856 6724
rect 384908 6712 384914 6724
rect 481726 6712 481732 6724
rect 384908 6684 481732 6712
rect 384908 6672 384914 6684
rect 481726 6672 481732 6684
rect 481784 6672 481790 6724
rect 130562 6604 130568 6656
rect 130620 6644 130626 6656
rect 274818 6644 274824 6656
rect 130620 6616 274824 6644
rect 130620 6604 130626 6616
rect 274818 6604 274824 6616
rect 274876 6604 274882 6656
rect 384758 6604 384764 6656
rect 384816 6644 384822 6656
rect 485222 6644 485228 6656
rect 384816 6616 485228 6644
rect 384816 6604 384822 6616
rect 485222 6604 485228 6616
rect 485280 6604 485286 6656
rect 69106 6536 69112 6588
rect 69164 6576 69170 6588
rect 255406 6576 255412 6588
rect 69164 6548 255412 6576
rect 69164 6536 69170 6548
rect 255406 6536 255412 6548
rect 255464 6536 255470 6588
rect 386322 6536 386328 6588
rect 386380 6576 386386 6588
rect 488810 6576 488816 6588
rect 386380 6548 488816 6576
rect 386380 6536 386386 6548
rect 488810 6536 488816 6548
rect 488868 6536 488874 6588
rect 65518 6468 65524 6520
rect 65576 6508 65582 6520
rect 254026 6508 254032 6520
rect 65576 6480 254032 6508
rect 65576 6468 65582 6480
rect 254026 6468 254032 6480
rect 254084 6468 254090 6520
rect 387702 6468 387708 6520
rect 387760 6508 387766 6520
rect 492306 6508 492312 6520
rect 387760 6480 492312 6508
rect 387760 6468 387766 6480
rect 492306 6468 492312 6480
rect 492364 6468 492370 6520
rect 62022 6400 62028 6452
rect 62080 6440 62086 6452
rect 254118 6440 254124 6452
rect 62080 6412 254124 6440
rect 62080 6400 62086 6412
rect 254118 6400 254124 6412
rect 254176 6400 254182 6452
rect 389082 6400 389088 6452
rect 389140 6440 389146 6452
rect 495894 6440 495900 6452
rect 389140 6412 495900 6440
rect 389140 6400 389146 6412
rect 495894 6400 495900 6412
rect 495952 6400 495958 6452
rect 58434 6332 58440 6384
rect 58492 6372 58498 6384
rect 252646 6372 252652 6384
rect 58492 6344 252652 6372
rect 58492 6332 58498 6344
rect 252646 6332 252652 6344
rect 252704 6332 252710 6384
rect 299658 6332 299664 6384
rect 299716 6372 299722 6384
rect 316678 6372 316684 6384
rect 299716 6344 316684 6372
rect 299716 6332 299722 6344
rect 316678 6332 316684 6344
rect 316736 6332 316742 6384
rect 390186 6332 390192 6384
rect 390244 6372 390250 6384
rect 499390 6372 499396 6384
rect 390244 6344 499396 6372
rect 390244 6332 390250 6344
rect 499390 6332 499396 6344
rect 499448 6332 499454 6384
rect 54938 6264 54944 6316
rect 54996 6304 55002 6316
rect 251358 6304 251364 6316
rect 54996 6276 251364 6304
rect 54996 6264 55002 6276
rect 251358 6264 251364 6276
rect 251416 6264 251422 6316
rect 259454 6264 259460 6316
rect 259512 6304 259518 6316
rect 295978 6304 295984 6316
rect 259512 6276 295984 6304
rect 259512 6264 259518 6276
rect 295978 6264 295984 6276
rect 296036 6264 296042 6316
rect 303154 6264 303160 6316
rect 303212 6304 303218 6316
rect 327718 6304 327724 6316
rect 303212 6276 327724 6304
rect 303212 6264 303218 6276
rect 327718 6264 327724 6276
rect 327776 6264 327782 6316
rect 390370 6264 390376 6316
rect 390428 6304 390434 6316
rect 502886 6304 502892 6316
rect 390428 6276 502892 6304
rect 390428 6264 390434 6276
rect 502886 6264 502892 6276
rect 502944 6264 502950 6316
rect 51350 6196 51356 6248
rect 51408 6236 51414 6248
rect 250070 6236 250076 6248
rect 51408 6208 250076 6236
rect 51408 6196 51414 6208
rect 250070 6196 250076 6208
rect 250128 6196 250134 6248
rect 268838 6196 268844 6248
rect 268896 6236 268902 6248
rect 317690 6236 317696 6248
rect 268896 6208 317696 6236
rect 268896 6196 268902 6208
rect 317690 6196 317696 6208
rect 317748 6196 317754 6248
rect 371878 6196 371884 6248
rect 371936 6236 371942 6248
rect 378870 6236 378876 6248
rect 371936 6208 378876 6236
rect 371936 6196 371942 6208
rect 378870 6196 378876 6208
rect 378928 6196 378934 6248
rect 391658 6196 391664 6248
rect 391716 6236 391722 6248
rect 506474 6236 506480 6248
rect 391716 6208 506480 6236
rect 391716 6196 391722 6208
rect 506474 6196 506480 6208
rect 506532 6196 506538 6248
rect 47854 6128 47860 6180
rect 47912 6168 47918 6180
rect 248506 6168 248512 6180
rect 47912 6140 248512 6168
rect 47912 6128 47918 6140
rect 248506 6128 248512 6140
rect 248564 6128 248570 6180
rect 257062 6128 257068 6180
rect 257120 6168 257126 6180
rect 313274 6168 313280 6180
rect 257120 6140 313280 6168
rect 257120 6128 257126 6140
rect 313274 6128 313280 6140
rect 313332 6128 313338 6180
rect 370498 6128 370504 6180
rect 370556 6168 370562 6180
rect 385954 6168 385960 6180
rect 370556 6140 385960 6168
rect 370556 6128 370562 6140
rect 385954 6128 385960 6140
rect 386012 6128 386018 6180
rect 393130 6128 393136 6180
rect 393188 6168 393194 6180
rect 510062 6168 510068 6180
rect 393188 6140 510068 6168
rect 393188 6128 393194 6140
rect 510062 6128 510068 6140
rect 510120 6128 510126 6180
rect 173158 6060 173164 6112
rect 173216 6100 173222 6112
rect 287146 6100 287152 6112
rect 173216 6072 287152 6100
rect 173216 6060 173222 6072
rect 287146 6060 287152 6072
rect 287204 6060 287210 6112
rect 382090 6060 382096 6112
rect 382148 6100 382154 6112
rect 473446 6100 473452 6112
rect 382148 6072 473452 6100
rect 382148 6060 382154 6072
rect 473446 6060 473452 6072
rect 473504 6060 473510 6112
rect 176654 5992 176660 6044
rect 176712 6032 176718 6044
rect 288618 6032 288624 6044
rect 176712 6004 288624 6032
rect 176712 5992 176718 6004
rect 288618 5992 288624 6004
rect 288676 5992 288682 6044
rect 380710 5992 380716 6044
rect 380768 6032 380774 6044
rect 469858 6032 469864 6044
rect 380768 6004 469864 6032
rect 380768 5992 380774 6004
rect 469858 5992 469864 6004
rect 469916 5992 469922 6044
rect 180242 5924 180248 5976
rect 180300 5964 180306 5976
rect 289998 5964 290004 5976
rect 180300 5936 290004 5964
rect 180300 5924 180306 5936
rect 289998 5924 290004 5936
rect 290056 5924 290062 5976
rect 379422 5924 379428 5976
rect 379480 5964 379486 5976
rect 466270 5964 466276 5976
rect 379480 5936 466276 5964
rect 379480 5924 379486 5936
rect 466270 5924 466276 5936
rect 466328 5924 466334 5976
rect 468478 5924 468484 5976
rect 468536 5964 468542 5976
rect 474550 5964 474556 5976
rect 468536 5936 474556 5964
rect 468536 5924 468542 5936
rect 474550 5924 474556 5936
rect 474608 5924 474614 5976
rect 183738 5856 183744 5908
rect 183796 5896 183802 5908
rect 291378 5896 291384 5908
rect 183796 5868 291384 5896
rect 183796 5856 183802 5868
rect 291378 5856 291384 5868
rect 291436 5856 291442 5908
rect 377950 5856 377956 5908
rect 378008 5896 378014 5908
rect 462774 5896 462780 5908
rect 378008 5868 462780 5896
rect 378008 5856 378014 5868
rect 462774 5856 462780 5868
rect 462832 5856 462838 5908
rect 187326 5788 187332 5840
rect 187384 5828 187390 5840
rect 292666 5828 292672 5840
rect 187384 5800 292672 5828
rect 187384 5788 187390 5800
rect 292666 5788 292672 5800
rect 292724 5788 292730 5840
rect 377858 5788 377864 5840
rect 377916 5828 377922 5840
rect 459186 5828 459192 5840
rect 377916 5800 459192 5828
rect 377916 5788 377922 5800
rect 459186 5788 459192 5800
rect 459244 5788 459250 5840
rect 190822 5720 190828 5772
rect 190880 5760 190886 5772
rect 292758 5760 292764 5772
rect 190880 5732 292764 5760
rect 190880 5720 190886 5732
rect 292758 5720 292764 5732
rect 292816 5720 292822 5772
rect 376662 5720 376668 5772
rect 376720 5760 376726 5772
rect 455690 5760 455696 5772
rect 376720 5732 455696 5760
rect 376720 5720 376726 5732
rect 455690 5720 455696 5732
rect 455748 5720 455754 5772
rect 194410 5652 194416 5704
rect 194468 5692 194474 5704
rect 294230 5692 294236 5704
rect 194468 5664 294236 5692
rect 194468 5652 194474 5664
rect 294230 5652 294236 5664
rect 294288 5652 294294 5704
rect 375190 5652 375196 5704
rect 375248 5692 375254 5704
rect 452102 5692 452108 5704
rect 375248 5664 452108 5692
rect 375248 5652 375254 5664
rect 452102 5652 452108 5664
rect 452160 5652 452166 5704
rect 363598 5516 363604 5568
rect 363656 5556 363662 5568
rect 367002 5556 367008 5568
rect 363656 5528 367008 5556
rect 363656 5516 363662 5528
rect 367002 5516 367008 5528
rect 367060 5516 367066 5568
rect 475378 5516 475384 5568
rect 475436 5556 475442 5568
rect 480530 5556 480536 5568
rect 475436 5528 480536 5556
rect 475436 5516 475442 5528
rect 480530 5516 480536 5528
rect 480588 5516 480594 5568
rect 486418 5516 486424 5568
rect 486476 5556 486482 5568
rect 487614 5556 487620 5568
rect 486476 5528 487620 5556
rect 486476 5516 486482 5528
rect 487614 5516 487620 5528
rect 487672 5516 487678 5568
rect 497458 5516 497464 5568
rect 497516 5556 497522 5568
rect 498194 5556 498200 5568
rect 497516 5528 498200 5556
rect 497516 5516 497522 5528
rect 498194 5516 498200 5528
rect 498252 5516 498258 5568
rect 504358 5516 504364 5568
rect 504416 5556 504422 5568
rect 505370 5556 505376 5568
rect 504416 5528 505376 5556
rect 504416 5516 504422 5528
rect 505370 5516 505376 5528
rect 505428 5516 505434 5568
rect 186130 5448 186136 5500
rect 186188 5488 186194 5500
rect 215938 5488 215944 5500
rect 186188 5460 215944 5488
rect 186188 5448 186194 5460
rect 215938 5448 215944 5460
rect 215996 5448 216002 5500
rect 218054 5448 218060 5500
rect 218112 5488 218118 5500
rect 302510 5488 302516 5500
rect 218112 5460 302516 5488
rect 218112 5448 218118 5460
rect 302510 5448 302516 5460
rect 302568 5448 302574 5500
rect 355870 5448 355876 5500
rect 355928 5488 355934 5500
rect 391842 5488 391848 5500
rect 355928 5460 391848 5488
rect 355928 5448 355934 5460
rect 391842 5448 391848 5460
rect 391900 5448 391906 5500
rect 402698 5448 402704 5500
rect 402756 5488 402762 5500
rect 540790 5488 540796 5500
rect 402756 5460 540796 5488
rect 402756 5448 402762 5460
rect 540790 5448 540796 5460
rect 540848 5448 540854 5500
rect 189718 5380 189724 5432
rect 189776 5420 189782 5432
rect 214282 5420 214288 5432
rect 189776 5392 214288 5420
rect 189776 5380 189782 5392
rect 214282 5380 214288 5392
rect 214340 5380 214346 5432
rect 214466 5380 214472 5432
rect 214524 5420 214530 5432
rect 301038 5420 301044 5432
rect 214524 5392 301044 5420
rect 214524 5380 214530 5392
rect 301038 5380 301044 5392
rect 301096 5380 301102 5432
rect 357250 5380 357256 5432
rect 357308 5420 357314 5432
rect 395246 5420 395252 5432
rect 357308 5392 395252 5420
rect 357308 5380 357314 5392
rect 395246 5380 395252 5392
rect 395304 5380 395310 5432
rect 404170 5380 404176 5432
rect 404228 5420 404234 5432
rect 544378 5420 544384 5432
rect 404228 5392 544384 5420
rect 404228 5380 404234 5392
rect 544378 5380 544384 5392
rect 544436 5380 544442 5432
rect 210970 5312 210976 5364
rect 211028 5352 211034 5364
rect 299750 5352 299756 5364
rect 211028 5324 299756 5352
rect 211028 5312 211034 5324
rect 299750 5312 299756 5324
rect 299808 5312 299814 5364
rect 358630 5312 358636 5364
rect 358688 5352 358694 5364
rect 400122 5352 400128 5364
rect 358688 5324 400128 5352
rect 358688 5312 358694 5324
rect 400122 5312 400128 5324
rect 400180 5312 400186 5364
rect 404078 5312 404084 5364
rect 404136 5352 404142 5364
rect 547874 5352 547880 5364
rect 404136 5324 547880 5352
rect 404136 5312 404142 5324
rect 547874 5312 547880 5324
rect 547932 5312 547938 5364
rect 136450 5244 136456 5296
rect 136508 5284 136514 5296
rect 204898 5284 204904 5296
rect 136508 5256 204904 5284
rect 136508 5244 136514 5256
rect 204898 5244 204904 5256
rect 204956 5244 204962 5296
rect 207382 5244 207388 5296
rect 207440 5284 207446 5296
rect 298278 5284 298284 5296
rect 207440 5256 298284 5284
rect 207440 5244 207446 5256
rect 298278 5244 298284 5256
rect 298336 5244 298342 5296
rect 358538 5244 358544 5296
rect 358596 5284 358602 5296
rect 398926 5284 398932 5296
rect 358596 5256 398932 5284
rect 358596 5244 358602 5256
rect 398926 5244 398932 5256
rect 398984 5244 398990 5296
rect 405550 5244 405556 5296
rect 405608 5284 405614 5296
rect 551462 5284 551468 5296
rect 405608 5256 551468 5284
rect 405608 5244 405614 5256
rect 551462 5244 551468 5256
rect 551520 5244 551526 5296
rect 203886 5176 203892 5228
rect 203944 5216 203950 5228
rect 296898 5216 296904 5228
rect 203944 5188 296904 5216
rect 203944 5176 203950 5188
rect 296898 5176 296904 5188
rect 296956 5176 296962 5228
rect 359918 5176 359924 5228
rect 359976 5216 359982 5228
rect 402514 5216 402520 5228
rect 359976 5188 402520 5216
rect 359976 5176 359982 5188
rect 402514 5176 402520 5188
rect 402572 5176 402578 5228
rect 406838 5176 406844 5228
rect 406896 5216 406902 5228
rect 554958 5216 554964 5228
rect 406896 5188 554964 5216
rect 406896 5176 406902 5188
rect 554958 5176 554964 5188
rect 555016 5176 555022 5228
rect 132954 5108 132960 5160
rect 133012 5148 133018 5160
rect 274726 5148 274732 5160
rect 133012 5120 274732 5148
rect 133012 5108 133018 5120
rect 274726 5108 274732 5120
rect 274784 5108 274790 5160
rect 278314 5108 278320 5160
rect 278372 5148 278378 5160
rect 320358 5148 320364 5160
rect 278372 5120 320364 5148
rect 278372 5108 278378 5120
rect 320358 5108 320364 5120
rect 320416 5108 320422 5160
rect 359826 5108 359832 5160
rect 359884 5148 359890 5160
rect 403618 5148 403624 5160
rect 359884 5120 403624 5148
rect 359884 5108 359890 5120
rect 403618 5108 403624 5120
rect 403676 5108 403682 5160
rect 408310 5108 408316 5160
rect 408368 5148 408374 5160
rect 558546 5148 558552 5160
rect 408368 5120 558552 5148
rect 408368 5108 408374 5120
rect 558546 5108 558552 5120
rect 558604 5108 558610 5160
rect 129366 5040 129372 5092
rect 129424 5080 129430 5092
rect 274634 5080 274640 5092
rect 129424 5052 274640 5080
rect 129424 5040 129430 5052
rect 274634 5040 274640 5052
rect 274692 5040 274698 5092
rect 274818 5040 274824 5092
rect 274876 5080 274882 5092
rect 318886 5080 318892 5092
rect 274876 5052 318892 5080
rect 274876 5040 274882 5052
rect 318886 5040 318892 5052
rect 318944 5040 318950 5092
rect 361298 5040 361304 5092
rect 361356 5080 361362 5092
rect 406010 5080 406016 5092
rect 361356 5052 406016 5080
rect 361356 5040 361362 5052
rect 406010 5040 406016 5052
rect 406068 5040 406074 5092
rect 409598 5040 409604 5092
rect 409656 5080 409662 5092
rect 562042 5080 562048 5092
rect 409656 5052 562048 5080
rect 409656 5040 409662 5052
rect 562042 5040 562048 5052
rect 562100 5040 562106 5092
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 236086 5012 236092 5024
rect 7708 4984 236092 5012
rect 7708 4972 7714 4984
rect 236086 4972 236092 4984
rect 236144 4972 236150 5024
rect 246390 4972 246396 5024
rect 246448 5012 246454 5024
rect 310514 5012 310520 5024
rect 246448 4984 310520 5012
rect 246448 4972 246454 4984
rect 310514 4972 310520 4984
rect 310572 4972 310578 5024
rect 361390 4972 361396 5024
rect 361448 5012 361454 5024
rect 407206 5012 407212 5024
rect 361448 4984 407212 5012
rect 361448 4972 361454 4984
rect 407206 4972 407212 4984
rect 407264 4972 407270 5024
rect 409690 4972 409696 5024
rect 409748 5012 409754 5024
rect 565630 5012 565636 5024
rect 409748 4984 565636 5012
rect 409748 4972 409754 4984
rect 565630 4972 565636 4984
rect 565688 4972 565694 5024
rect 2866 4904 2872 4956
rect 2924 4944 2930 4956
rect 234706 4944 234712 4956
rect 2924 4916 234712 4944
rect 2924 4904 2930 4916
rect 234706 4904 234712 4916
rect 234764 4904 234770 4956
rect 242894 4904 242900 4956
rect 242952 4944 242958 4956
rect 309134 4944 309140 4956
rect 242952 4916 309140 4944
rect 242952 4904 242958 4916
rect 309134 4904 309140 4916
rect 309192 4904 309198 4956
rect 362678 4904 362684 4956
rect 362736 4944 362742 4956
rect 410794 4944 410800 4956
rect 362736 4916 410800 4944
rect 362736 4904 362742 4916
rect 410794 4904 410800 4916
rect 410852 4904 410858 4956
rect 411070 4904 411076 4956
rect 411128 4944 411134 4956
rect 569126 4944 569132 4956
rect 411128 4916 569132 4944
rect 411128 4904 411134 4916
rect 569126 4904 569132 4916
rect 569184 4904 569190 4956
rect 1670 4836 1676 4888
rect 1728 4876 1734 4888
rect 234798 4876 234804 4888
rect 1728 4848 234804 4876
rect 1728 4836 1734 4848
rect 234798 4836 234804 4848
rect 234856 4836 234862 4888
rect 239306 4836 239312 4888
rect 239364 4876 239370 4888
rect 307754 4876 307760 4888
rect 239364 4848 307760 4876
rect 239364 4836 239370 4848
rect 307754 4836 307760 4848
rect 307812 4836 307818 4888
rect 361206 4836 361212 4888
rect 361264 4876 361270 4888
rect 409598 4876 409604 4888
rect 361264 4848 409604 4876
rect 361264 4836 361270 4848
rect 409598 4836 409604 4848
rect 409656 4836 409662 4888
rect 412358 4836 412364 4888
rect 412416 4876 412422 4888
rect 572714 4876 572720 4888
rect 412416 4848 572720 4876
rect 412416 4836 412422 4848
rect 572714 4836 572720 4848
rect 572772 4836 572778 4888
rect 566 4768 572 4820
rect 624 4808 630 4820
rect 234890 4808 234896 4820
rect 624 4780 234896 4808
rect 624 4768 630 4780
rect 234890 4768 234896 4780
rect 234948 4768 234954 4820
rect 235810 4768 235816 4820
rect 235868 4808 235874 4820
rect 306374 4808 306380 4820
rect 235868 4780 306380 4808
rect 235868 4768 235874 4780
rect 306374 4768 306380 4780
rect 306432 4768 306438 4820
rect 362770 4768 362776 4820
rect 362828 4808 362834 4820
rect 413094 4808 413100 4820
rect 362828 4780 413100 4808
rect 362828 4768 362834 4780
rect 413094 4768 413100 4780
rect 413152 4768 413158 4820
rect 413830 4768 413836 4820
rect 413888 4808 413894 4820
rect 576302 4808 576308 4820
rect 413888 4780 576308 4808
rect 413888 4768 413894 4780
rect 576302 4768 576308 4780
rect 576360 4768 576366 4820
rect 193214 4700 193220 4752
rect 193272 4740 193278 4752
rect 220078 4740 220084 4752
rect 193272 4712 220084 4740
rect 193272 4700 193278 4712
rect 220078 4700 220084 4712
rect 220136 4700 220142 4752
rect 221550 4700 221556 4752
rect 221608 4740 221614 4752
rect 302326 4740 302332 4752
rect 221608 4712 302332 4740
rect 221608 4700 221614 4712
rect 302326 4700 302332 4712
rect 302384 4700 302390 4752
rect 355778 4700 355784 4752
rect 355836 4740 355842 4752
rect 388254 4740 388260 4752
rect 355836 4712 388260 4740
rect 355836 4700 355842 4712
rect 388254 4700 388260 4712
rect 388312 4700 388318 4752
rect 401318 4700 401324 4752
rect 401376 4740 401382 4752
rect 537202 4740 537208 4752
rect 401376 4712 537208 4740
rect 401376 4700 401382 4712
rect 537202 4700 537208 4712
rect 537260 4700 537266 4752
rect 171962 4632 171968 4684
rect 172020 4672 172026 4684
rect 222838 4672 222844 4684
rect 172020 4644 222844 4672
rect 172020 4632 172026 4644
rect 222838 4632 222844 4644
rect 222896 4632 222902 4684
rect 225138 4632 225144 4684
rect 225196 4672 225202 4684
rect 303798 4672 303804 4684
rect 225196 4644 303804 4672
rect 225196 4632 225202 4644
rect 303798 4632 303804 4644
rect 303856 4632 303862 4684
rect 354490 4632 354496 4684
rect 354548 4672 354554 4684
rect 384758 4672 384764 4684
rect 354548 4644 384764 4672
rect 354548 4632 354554 4644
rect 384758 4632 384764 4644
rect 384816 4632 384822 4684
rect 399846 4632 399852 4684
rect 399904 4672 399910 4684
rect 533706 4672 533712 4684
rect 399904 4644 533712 4672
rect 399904 4632 399910 4644
rect 533706 4632 533712 4644
rect 533764 4632 533770 4684
rect 228726 4564 228732 4616
rect 228784 4604 228790 4616
rect 304994 4604 305000 4616
rect 228784 4576 305000 4604
rect 228784 4564 228790 4576
rect 304994 4564 305000 4576
rect 305052 4564 305058 4616
rect 353110 4564 353116 4616
rect 353168 4604 353174 4616
rect 381170 4604 381176 4616
rect 353168 4576 381176 4604
rect 353168 4564 353174 4576
rect 381170 4564 381176 4576
rect 381228 4564 381234 4616
rect 398650 4564 398656 4616
rect 398708 4604 398714 4616
rect 530118 4604 530124 4616
rect 398708 4576 530124 4604
rect 398708 4564 398714 4576
rect 530118 4564 530124 4576
rect 530176 4564 530182 4616
rect 232222 4496 232228 4548
rect 232280 4536 232286 4548
rect 306466 4536 306472 4548
rect 232280 4508 306472 4536
rect 232280 4496 232286 4508
rect 306466 4496 306472 4508
rect 306524 4496 306530 4548
rect 351730 4496 351736 4548
rect 351788 4536 351794 4548
rect 377674 4536 377680 4548
rect 351788 4508 377680 4536
rect 351788 4496 351794 4508
rect 377674 4496 377680 4508
rect 377732 4496 377738 4548
rect 398558 4496 398564 4548
rect 398616 4536 398622 4548
rect 526622 4536 526628 4548
rect 398616 4508 526628 4536
rect 398616 4496 398622 4508
rect 526622 4496 526628 4508
rect 526680 4496 526686 4548
rect 281902 4428 281908 4480
rect 281960 4468 281966 4480
rect 321738 4468 321744 4480
rect 281960 4440 321744 4468
rect 281960 4428 281966 4440
rect 321738 4428 321744 4440
rect 321796 4428 321802 4480
rect 350258 4428 350264 4480
rect 350316 4468 350322 4480
rect 374086 4468 374092 4480
rect 350316 4440 374092 4468
rect 350316 4428 350322 4440
rect 374086 4428 374092 4440
rect 374144 4428 374150 4480
rect 397086 4428 397092 4480
rect 397144 4468 397150 4480
rect 523034 4468 523040 4480
rect 397144 4440 523040 4468
rect 397144 4428 397150 4440
rect 523034 4428 523040 4440
rect 523092 4428 523098 4480
rect 285398 4360 285404 4412
rect 285456 4400 285462 4412
rect 323026 4400 323032 4412
rect 285456 4372 323032 4400
rect 285456 4360 285462 4372
rect 323026 4360 323032 4372
rect 323084 4360 323090 4412
rect 395798 4360 395804 4412
rect 395856 4400 395862 4412
rect 519538 4400 519544 4412
rect 395856 4372 519544 4400
rect 395856 4360 395862 4372
rect 519538 4360 519544 4372
rect 519596 4360 519602 4412
rect 288986 4292 288992 4344
rect 289044 4332 289050 4344
rect 323118 4332 323124 4344
rect 289044 4304 323124 4332
rect 289044 4292 289050 4304
rect 323118 4292 323124 4304
rect 323176 4292 323182 4344
rect 394418 4292 394424 4344
rect 394476 4332 394482 4344
rect 515950 4332 515956 4344
rect 394476 4304 515956 4332
rect 394476 4292 394482 4304
rect 515950 4292 515956 4304
rect 516008 4292 516014 4344
rect 200298 4224 200304 4276
rect 200356 4264 200362 4276
rect 208946 4264 208952 4276
rect 200356 4236 208952 4264
rect 200356 4224 200362 4236
rect 208946 4224 208952 4236
rect 209004 4224 209010 4276
rect 292574 4224 292580 4276
rect 292632 4264 292638 4276
rect 324590 4264 324596 4276
rect 292632 4236 324596 4264
rect 292632 4224 292638 4236
rect 324590 4224 324596 4236
rect 324648 4224 324654 4276
rect 392946 4224 392952 4276
rect 393004 4264 393010 4276
rect 512454 4264 512460 4276
rect 393004 4236 512460 4264
rect 393004 4224 393010 4236
rect 512454 4224 512460 4236
rect 512512 4224 512518 4276
rect 84028 4168 84516 4196
rect 11146 4088 11152 4140
rect 11204 4128 11210 4140
rect 18598 4128 18604 4140
rect 11204 4100 18604 4128
rect 11204 4088 11210 4100
rect 18598 4088 18604 4100
rect 18656 4088 18662 4140
rect 34790 4088 34796 4140
rect 34848 4128 34854 4140
rect 36538 4128 36544 4140
rect 34848 4100 36544 4128
rect 34848 4088 34854 4100
rect 36538 4088 36544 4100
rect 36596 4088 36602 4140
rect 78490 4088 78496 4140
rect 78548 4128 78554 4140
rect 84028 4128 84056 4168
rect 78548 4100 84056 4128
rect 78548 4088 78554 4100
rect 82078 4020 82084 4072
rect 82136 4060 82142 4072
rect 84289 4063 84347 4069
rect 84289 4060 84301 4063
rect 82136 4032 84301 4060
rect 82136 4020 82142 4032
rect 84289 4029 84301 4032
rect 84335 4029 84347 4063
rect 84488 4060 84516 4168
rect 143534 4156 143540 4208
rect 143592 4196 143598 4208
rect 144822 4196 144828 4208
rect 143592 4168 144828 4196
rect 143592 4156 143598 4168
rect 144822 4156 144828 4168
rect 144880 4156 144886 4208
rect 168374 4156 168380 4208
rect 168432 4196 168438 4208
rect 169662 4196 169668 4208
rect 168432 4168 169668 4196
rect 168432 4156 168438 4168
rect 169662 4156 169668 4168
rect 169720 4156 169726 4208
rect 201494 4156 201500 4208
rect 201552 4196 201558 4208
rect 202782 4196 202788 4208
rect 201552 4168 202788 4196
rect 201552 4156 201558 4168
rect 202782 4156 202788 4168
rect 202840 4156 202846 4208
rect 226334 4156 226340 4208
rect 226392 4196 226398 4208
rect 227622 4196 227628 4208
rect 226392 4168 227628 4196
rect 226392 4156 226398 4168
rect 227622 4156 227628 4168
rect 227680 4156 227686 4208
rect 388438 4156 388444 4208
rect 388496 4196 388502 4208
rect 389450 4196 389456 4208
rect 388496 4168 389456 4196
rect 388496 4156 388502 4168
rect 389450 4156 389456 4168
rect 389508 4156 389514 4208
rect 395338 4156 395344 4208
rect 395396 4196 395402 4208
rect 396534 4196 396540 4208
rect 395396 4168 396540 4196
rect 395396 4156 395402 4168
rect 396534 4156 396540 4168
rect 396592 4156 396598 4208
rect 84565 4131 84623 4137
rect 84565 4097 84577 4131
rect 84611 4128 84623 4131
rect 259730 4128 259736 4140
rect 84611 4100 259736 4128
rect 84611 4097 84623 4100
rect 84565 4091 84623 4097
rect 259730 4088 259736 4100
rect 259788 4088 259794 4140
rect 309042 4088 309048 4140
rect 309100 4128 309106 4140
rect 330110 4128 330116 4140
rect 309100 4100 330116 4128
rect 309100 4088 309106 4100
rect 330110 4088 330116 4100
rect 330168 4088 330174 4140
rect 332686 4088 332692 4140
rect 332744 4128 332750 4140
rect 335998 4128 336004 4140
rect 332744 4100 336004 4128
rect 332744 4088 332750 4100
rect 335998 4088 336004 4100
rect 336056 4088 336062 4140
rect 343450 4088 343456 4140
rect 343508 4128 343514 4140
rect 350442 4128 350448 4140
rect 343508 4100 350448 4128
rect 343508 4088 343514 4100
rect 350442 4088 350448 4100
rect 350500 4088 350506 4140
rect 351822 4088 351828 4140
rect 351880 4128 351886 4140
rect 375282 4128 375288 4140
rect 351880 4100 375288 4128
rect 351880 4088 351886 4100
rect 375282 4088 375288 4100
rect 375340 4088 375346 4140
rect 402606 4088 402612 4140
rect 402664 4128 402670 4140
rect 534997 4131 535055 4137
rect 534997 4128 535009 4131
rect 402664 4100 535009 4128
rect 402664 4088 402670 4100
rect 534997 4097 535009 4100
rect 535043 4097 535055 4131
rect 534997 4091 535055 4097
rect 258166 4060 258172 4072
rect 84488 4032 258172 4060
rect 84289 4023 84347 4029
rect 258166 4020 258172 4032
rect 258224 4020 258230 4072
rect 307938 4020 307944 4072
rect 307996 4060 308002 4072
rect 330018 4060 330024 4072
rect 307996 4032 330024 4060
rect 307996 4020 308002 4032
rect 330018 4020 330024 4032
rect 330076 4020 330082 4072
rect 343542 4020 343548 4072
rect 343600 4060 343606 4072
rect 348050 4060 348056 4072
rect 343600 4032 348056 4060
rect 343600 4020 343606 4032
rect 348050 4020 348056 4032
rect 348108 4020 348114 4072
rect 350350 4020 350356 4072
rect 350408 4060 350414 4072
rect 372890 4060 372896 4072
rect 350408 4032 372896 4060
rect 350408 4020 350414 4032
rect 372890 4020 372896 4032
rect 372948 4020 372954 4072
rect 402790 4020 402796 4072
rect 402848 4060 402854 4072
rect 543182 4060 543188 4072
rect 402848 4032 543188 4060
rect 402848 4020 402854 4032
rect 543182 4020 543188 4032
rect 543240 4020 543246 4072
rect 43070 3952 43076 4004
rect 43128 3992 43134 4004
rect 51718 3992 51724 4004
rect 43128 3964 51724 3992
rect 43128 3952 43134 3964
rect 51718 3952 51724 3964
rect 51776 3952 51782 4004
rect 53650 3952 53656 4004
rect 53708 3992 53714 4004
rect 57238 3992 57244 4004
rect 53708 3964 57244 3992
rect 53708 3952 53714 3964
rect 57238 3952 57244 3964
rect 57296 3952 57302 4004
rect 74994 3952 75000 4004
rect 75052 3992 75058 4004
rect 258074 3992 258080 4004
rect 75052 3964 258080 3992
rect 75052 3952 75058 3964
rect 258074 3952 258080 3964
rect 258132 3952 258138 4004
rect 305546 3952 305552 4004
rect 305604 3992 305610 4004
rect 328546 3992 328552 4004
rect 305604 3964 328552 3992
rect 305604 3952 305610 3964
rect 328546 3952 328552 3964
rect 328604 3952 328610 4004
rect 329190 3952 329196 4004
rect 329248 3992 329254 4004
rect 335446 3992 335452 4004
rect 329248 3964 335452 3992
rect 329248 3952 329254 3964
rect 335446 3952 335452 3964
rect 335504 3952 335510 4004
rect 343358 3952 343364 4004
rect 343416 3992 343422 4004
rect 349246 3992 349252 4004
rect 343416 3964 349252 3992
rect 343416 3952 343422 3964
rect 349246 3952 349252 3964
rect 349304 3952 349310 4004
rect 353202 3952 353208 4004
rect 353260 3992 353266 4004
rect 379974 3992 379980 4004
rect 353260 3964 379980 3992
rect 353260 3952 353266 3964
rect 379974 3952 379980 3964
rect 380032 3952 380038 4004
rect 404262 3952 404268 4004
rect 404320 3992 404326 4004
rect 546678 3992 546684 4004
rect 404320 3964 546684 3992
rect 404320 3952 404326 3964
rect 546678 3952 546684 3964
rect 546736 3952 546742 4004
rect 38378 3884 38384 3936
rect 38436 3924 38442 3936
rect 47578 3924 47584 3936
rect 38436 3896 47584 3924
rect 38436 3884 38442 3896
rect 47578 3884 47584 3896
rect 47636 3884 47642 3936
rect 50154 3884 50160 3936
rect 50212 3924 50218 3936
rect 68278 3924 68284 3936
rect 50212 3896 68284 3924
rect 50212 3884 50218 3896
rect 68278 3884 68284 3896
rect 68336 3884 68342 3936
rect 71498 3884 71504 3936
rect 71556 3924 71562 3936
rect 256694 3924 256700 3936
rect 71556 3896 256700 3924
rect 71556 3884 71562 3896
rect 256694 3884 256700 3896
rect 256752 3884 256758 3936
rect 301958 3884 301964 3936
rect 302016 3924 302022 3936
rect 320729 3927 320787 3933
rect 320729 3924 320741 3927
rect 302016 3896 320741 3924
rect 302016 3884 302022 3896
rect 320729 3893 320741 3896
rect 320775 3893 320787 3927
rect 325786 3924 325792 3936
rect 320729 3887 320787 3893
rect 320836 3896 325792 3924
rect 5258 3816 5264 3868
rect 5316 3856 5322 3868
rect 7558 3856 7564 3868
rect 5316 3828 7564 3856
rect 5316 3816 5322 3828
rect 7558 3816 7564 3828
rect 7616 3816 7622 3868
rect 41874 3816 41880 3868
rect 41932 3856 41938 3868
rect 54478 3856 54484 3868
rect 41932 3828 54484 3856
rect 41932 3816 41938 3828
rect 54478 3816 54484 3828
rect 54536 3816 54542 3868
rect 67910 3816 67916 3868
rect 67968 3856 67974 3868
rect 255314 3856 255320 3868
rect 67968 3828 255320 3856
rect 67968 3816 67974 3828
rect 255314 3816 255320 3828
rect 255372 3816 255378 3868
rect 297266 3816 297272 3868
rect 297324 3856 297330 3868
rect 320836 3856 320864 3896
rect 325786 3884 325792 3896
rect 325844 3884 325850 3936
rect 334250 3924 334256 3936
rect 326356 3896 334256 3924
rect 297324 3828 320864 3856
rect 297324 3816 297330 3828
rect 320910 3816 320916 3868
rect 320968 3856 320974 3868
rect 326249 3859 326307 3865
rect 326249 3856 326261 3859
rect 320968 3828 326261 3856
rect 320968 3816 320974 3828
rect 326249 3825 326261 3828
rect 326295 3825 326307 3859
rect 326249 3819 326307 3825
rect 35986 3748 35992 3800
rect 36044 3788 36050 3800
rect 50338 3788 50344 3800
rect 36044 3760 50344 3788
rect 36044 3748 36050 3760
rect 50338 3748 50344 3760
rect 50396 3748 50402 3800
rect 64322 3748 64328 3800
rect 64380 3788 64386 3800
rect 253934 3788 253940 3800
rect 64380 3760 253940 3788
rect 64380 3748 64386 3760
rect 253934 3748 253940 3760
rect 253992 3748 253998 3800
rect 293678 3748 293684 3800
rect 293736 3788 293742 3800
rect 324314 3788 324320 3800
rect 293736 3760 324320 3788
rect 293736 3748 293742 3760
rect 324314 3748 324320 3760
rect 324372 3748 324378 3800
rect 324406 3748 324412 3800
rect 324464 3788 324470 3800
rect 326356 3788 326384 3896
rect 334250 3884 334256 3896
rect 334308 3884 334314 3936
rect 344278 3884 344284 3936
rect 344336 3924 344342 3936
rect 351638 3924 351644 3936
rect 344336 3896 351644 3924
rect 344336 3884 344342 3896
rect 351638 3884 351644 3896
rect 351696 3884 351702 3936
rect 354582 3884 354588 3936
rect 354640 3924 354646 3936
rect 387150 3924 387156 3936
rect 354640 3896 387156 3924
rect 354640 3884 354646 3896
rect 387150 3884 387156 3896
rect 387208 3884 387214 3936
rect 405642 3884 405648 3936
rect 405700 3924 405706 3936
rect 550266 3924 550272 3936
rect 405700 3896 550272 3924
rect 405700 3884 405706 3896
rect 550266 3884 550272 3896
rect 550324 3884 550330 3936
rect 326433 3859 326491 3865
rect 326433 3825 326445 3859
rect 326479 3856 326491 3859
rect 329098 3856 329104 3868
rect 326479 3828 329104 3856
rect 326479 3825 326491 3828
rect 326433 3819 326491 3825
rect 329098 3816 329104 3828
rect 329156 3816 329162 3868
rect 333882 3816 333888 3868
rect 333940 3856 333946 3868
rect 336918 3856 336924 3868
rect 333940 3828 336924 3856
rect 333940 3816 333946 3828
rect 336918 3816 336924 3828
rect 336976 3816 336982 3868
rect 345750 3816 345756 3868
rect 345808 3856 345814 3868
rect 356330 3856 356336 3868
rect 345808 3828 356336 3856
rect 345808 3816 345814 3828
rect 356330 3816 356336 3828
rect 356388 3816 356394 3868
rect 357342 3816 357348 3868
rect 357400 3856 357406 3868
rect 363785 3859 363843 3865
rect 357400 3828 363736 3856
rect 357400 3816 357406 3828
rect 327258 3788 327264 3800
rect 324464 3760 326384 3788
rect 326448 3760 327264 3788
rect 324464 3748 324470 3760
rect 23014 3680 23020 3732
rect 23072 3720 23078 3732
rect 39298 3720 39304 3732
rect 23072 3692 39304 3720
rect 23072 3680 23078 3692
rect 39298 3680 39304 3692
rect 39356 3680 39362 3732
rect 43438 3720 43444 3732
rect 39500 3692 43444 3720
rect 20622 3612 20628 3664
rect 20680 3652 20686 3664
rect 39500 3652 39528 3692
rect 43438 3680 43444 3692
rect 43496 3680 43502 3732
rect 45370 3680 45376 3732
rect 45428 3720 45434 3732
rect 58618 3720 58624 3732
rect 45428 3692 58624 3720
rect 45428 3680 45434 3692
rect 58618 3680 58624 3692
rect 58676 3680 58682 3732
rect 60826 3680 60832 3732
rect 60884 3720 60890 3732
rect 252830 3720 252836 3732
rect 60884 3692 252836 3720
rect 60884 3680 60890 3692
rect 252830 3680 252836 3692
rect 252888 3680 252894 3732
rect 291378 3680 291384 3732
rect 291436 3720 291442 3732
rect 320269 3723 320327 3729
rect 320269 3720 320281 3723
rect 291436 3692 320281 3720
rect 291436 3680 291442 3692
rect 320269 3689 320281 3692
rect 320315 3689 320327 3723
rect 320269 3683 320327 3689
rect 320729 3723 320787 3729
rect 320729 3689 320741 3723
rect 320775 3720 320787 3723
rect 326448 3720 326476 3760
rect 327258 3748 327264 3760
rect 327316 3748 327322 3800
rect 331214 3748 331220 3800
rect 331272 3788 331278 3800
rect 331490 3788 331496 3800
rect 331272 3760 331496 3788
rect 331272 3748 331278 3760
rect 331490 3748 331496 3760
rect 331548 3748 331554 3800
rect 346302 3748 346308 3800
rect 346360 3788 346366 3800
rect 346360 3760 354352 3788
rect 346360 3748 346366 3760
rect 320775 3692 326476 3720
rect 320775 3689 320787 3692
rect 320729 3683 320787 3689
rect 326798 3680 326804 3732
rect 326856 3720 326862 3732
rect 335630 3720 335636 3732
rect 326856 3692 335636 3720
rect 326856 3680 326862 3692
rect 335630 3680 335636 3692
rect 335688 3680 335694 3732
rect 347590 3680 347596 3732
rect 347648 3720 347654 3732
rect 354217 3723 354275 3729
rect 354217 3720 354229 3723
rect 347648 3692 354229 3720
rect 347648 3680 347654 3692
rect 354217 3689 354229 3692
rect 354263 3689 354275 3723
rect 354217 3683 354275 3689
rect 20680 3624 39528 3652
rect 20680 3612 20686 3624
rect 39574 3612 39580 3664
rect 39632 3652 39638 3664
rect 53929 3655 53987 3661
rect 39632 3624 53880 3652
rect 39632 3612 39638 3624
rect 18230 3544 18236 3596
rect 18288 3584 18294 3596
rect 18288 3556 26234 3584
rect 18288 3544 18294 3556
rect 26206 3516 26234 3556
rect 28902 3544 28908 3596
rect 28960 3584 28966 3596
rect 35158 3584 35164 3596
rect 28960 3556 35164 3584
rect 28960 3544 28966 3556
rect 35158 3544 35164 3556
rect 35216 3544 35222 3596
rect 40678 3544 40684 3596
rect 40736 3584 40742 3596
rect 41322 3584 41328 3596
rect 40736 3556 41328 3584
rect 40736 3544 40742 3556
rect 41322 3544 41328 3556
rect 41380 3544 41386 3596
rect 48958 3544 48964 3596
rect 49016 3584 49022 3596
rect 49602 3584 49608 3596
rect 49016 3556 49608 3584
rect 49016 3544 49022 3556
rect 49602 3544 49608 3556
rect 49660 3544 49666 3596
rect 52546 3544 52552 3596
rect 52604 3584 52610 3596
rect 53742 3584 53748 3596
rect 52604 3556 53748 3584
rect 52604 3544 52610 3556
rect 53742 3544 53748 3556
rect 53800 3544 53806 3596
rect 53852 3584 53880 3624
rect 53929 3621 53941 3655
rect 53975 3652 53987 3655
rect 248690 3652 248696 3664
rect 53975 3624 248696 3652
rect 53975 3621 53987 3624
rect 53929 3615 53987 3621
rect 248690 3612 248696 3624
rect 248748 3612 248754 3664
rect 286594 3612 286600 3664
rect 286652 3652 286658 3664
rect 323210 3652 323216 3664
rect 286652 3624 323216 3652
rect 286652 3612 286658 3624
rect 323210 3612 323216 3624
rect 323268 3612 323274 3664
rect 324222 3652 324228 3664
rect 323320 3624 324228 3652
rect 247218 3584 247224 3596
rect 53852 3556 247224 3584
rect 247218 3544 247224 3556
rect 247276 3544 247282 3596
rect 279510 3544 279516 3596
rect 279568 3584 279574 3596
rect 279568 3556 281580 3584
rect 279568 3544 279574 3556
rect 32306 3516 32312 3528
rect 26206 3488 32312 3516
rect 32306 3476 32312 3488
rect 32364 3476 32370 3528
rect 32398 3476 32404 3528
rect 32456 3516 32462 3528
rect 244458 3516 244464 3528
rect 32456 3488 244464 3516
rect 32456 3476 32462 3488
rect 244458 3476 244464 3488
rect 244516 3476 244522 3528
rect 249978 3476 249984 3528
rect 250036 3516 250042 3528
rect 251082 3516 251088 3528
rect 250036 3488 251088 3516
rect 250036 3476 250042 3488
rect 251082 3476 251088 3488
rect 251140 3476 251146 3528
rect 255866 3476 255872 3528
rect 255924 3516 255930 3528
rect 256602 3516 256608 3528
rect 255924 3488 256608 3516
rect 255924 3476 255930 3488
rect 256602 3476 256608 3488
rect 256660 3476 256666 3528
rect 262950 3476 262956 3528
rect 263008 3516 263014 3528
rect 263502 3516 263508 3528
rect 263008 3488 263508 3516
rect 263008 3476 263014 3488
rect 263502 3476 263508 3488
rect 263560 3476 263566 3528
rect 264146 3476 264152 3528
rect 264204 3516 264210 3528
rect 264882 3516 264888 3528
rect 264204 3488 264888 3516
rect 264204 3476 264210 3488
rect 264882 3476 264888 3488
rect 264940 3476 264946 3528
rect 266538 3476 266544 3528
rect 266596 3516 266602 3528
rect 267642 3516 267648 3528
rect 266596 3488 267648 3516
rect 266596 3476 266602 3488
rect 267642 3476 267648 3488
rect 267700 3476 267706 3528
rect 267734 3476 267740 3528
rect 267792 3516 267798 3528
rect 269022 3516 269028 3528
rect 267792 3488 269028 3516
rect 267792 3476 267798 3488
rect 269022 3476 269028 3488
rect 269080 3476 269086 3528
rect 271230 3476 271236 3528
rect 271288 3516 271294 3528
rect 271782 3516 271788 3528
rect 271288 3488 271788 3516
rect 271288 3476 271294 3488
rect 271782 3476 271788 3488
rect 271840 3476 271846 3528
rect 273622 3476 273628 3528
rect 273680 3516 273686 3528
rect 274542 3516 274548 3528
rect 273680 3488 274548 3516
rect 273680 3476 273686 3488
rect 274542 3476 274548 3488
rect 274600 3476 274606 3528
rect 280706 3476 280712 3528
rect 280764 3516 280770 3528
rect 281442 3516 281448 3528
rect 280764 3488 281448 3516
rect 280764 3476 280770 3488
rect 281442 3476 281448 3488
rect 281500 3476 281506 3528
rect 281552 3516 281580 3556
rect 284294 3544 284300 3596
rect 284352 3584 284358 3596
rect 321830 3584 321836 3596
rect 284352 3556 321836 3584
rect 284352 3544 284358 3556
rect 321830 3544 321836 3556
rect 321888 3544 321894 3596
rect 323320 3584 323348 3624
rect 324222 3612 324228 3624
rect 324280 3612 324286 3664
rect 325602 3612 325608 3664
rect 325660 3652 325666 3664
rect 335538 3652 335544 3664
rect 325660 3624 335544 3652
rect 325660 3612 325666 3624
rect 335538 3612 335544 3624
rect 335596 3612 335602 3664
rect 347130 3612 347136 3664
rect 347188 3652 347194 3664
rect 354324 3652 354352 3760
rect 358722 3748 358728 3800
rect 358780 3788 358786 3800
rect 363708 3788 363736 3828
rect 363785 3825 363797 3859
rect 363831 3856 363843 3859
rect 390646 3856 390652 3868
rect 363831 3828 390652 3856
rect 363831 3825 363843 3828
rect 363785 3819 363843 3825
rect 390646 3816 390652 3828
rect 390704 3816 390710 3868
rect 407022 3816 407028 3868
rect 407080 3856 407086 3868
rect 553762 3856 553768 3868
rect 407080 3828 553768 3856
rect 407080 3816 407086 3828
rect 553762 3816 553768 3828
rect 553820 3816 553826 3868
rect 394234 3788 394240 3800
rect 358780 3760 363644 3788
rect 363708 3760 394240 3788
rect 358780 3748 358786 3760
rect 358078 3680 358084 3732
rect 358136 3720 358142 3732
rect 363506 3720 363512 3732
rect 358136 3692 363512 3720
rect 358136 3680 358142 3692
rect 363506 3680 363512 3692
rect 363564 3680 363570 3732
rect 363616 3720 363644 3760
rect 394234 3748 394240 3760
rect 394292 3748 394298 3800
rect 406930 3748 406936 3800
rect 406988 3788 406994 3800
rect 557350 3788 557356 3800
rect 406988 3760 557356 3788
rect 406988 3748 406994 3760
rect 557350 3748 557356 3760
rect 557408 3748 557414 3800
rect 397730 3720 397736 3732
rect 363616 3692 397736 3720
rect 397730 3680 397736 3692
rect 397788 3680 397794 3732
rect 408402 3680 408408 3732
rect 408460 3720 408466 3732
rect 560846 3720 560852 3732
rect 408460 3692 560852 3720
rect 408460 3680 408466 3692
rect 560846 3680 560852 3692
rect 560904 3680 560910 3732
rect 358722 3652 358728 3664
rect 347188 3624 353064 3652
rect 354324 3624 358728 3652
rect 347188 3612 347194 3624
rect 321940 3556 323348 3584
rect 320174 3516 320180 3528
rect 281552 3488 320180 3516
rect 320174 3476 320180 3488
rect 320232 3476 320238 3528
rect 320269 3519 320327 3525
rect 320269 3485 320281 3519
rect 320315 3516 320327 3519
rect 321940 3516 321968 3556
rect 323394 3544 323400 3596
rect 323452 3584 323458 3596
rect 334066 3584 334072 3596
rect 323452 3556 334072 3584
rect 323452 3544 323458 3556
rect 334066 3544 334072 3556
rect 334124 3544 334130 3596
rect 342070 3544 342076 3596
rect 342128 3584 342134 3596
rect 346946 3584 346952 3596
rect 342128 3556 346952 3584
rect 342128 3544 342134 3556
rect 346946 3544 346952 3556
rect 347004 3544 347010 3596
rect 347682 3544 347688 3596
rect 347740 3584 347746 3596
rect 353036 3584 353064 3624
rect 358722 3612 358728 3624
rect 358780 3612 358786 3664
rect 360010 3612 360016 3664
rect 360068 3652 360074 3664
rect 401318 3652 401324 3664
rect 360068 3624 401324 3652
rect 360068 3612 360074 3624
rect 401318 3612 401324 3624
rect 401376 3612 401382 3664
rect 409782 3612 409788 3664
rect 409840 3652 409846 3664
rect 564434 3652 564440 3664
rect 409840 3624 564440 3652
rect 409840 3612 409846 3624
rect 564434 3612 564440 3624
rect 564492 3612 564498 3664
rect 359918 3584 359924 3596
rect 347740 3556 352972 3584
rect 353036 3556 359924 3584
rect 347740 3544 347746 3556
rect 320315 3488 321968 3516
rect 320315 3485 320327 3488
rect 320269 3479 320327 3485
rect 322106 3476 322112 3528
rect 322164 3516 322170 3528
rect 329929 3519 329987 3525
rect 329929 3516 329941 3519
rect 322164 3488 329941 3516
rect 322164 3476 322170 3488
rect 329929 3485 329941 3488
rect 329975 3485 329987 3519
rect 329929 3479 329987 3485
rect 331582 3476 331588 3528
rect 331640 3516 331646 3528
rect 332502 3516 332508 3528
rect 331640 3488 332508 3516
rect 331640 3476 331646 3488
rect 332502 3476 332508 3488
rect 332560 3476 332566 3528
rect 336274 3476 336280 3528
rect 336332 3516 336338 3528
rect 338114 3516 338120 3528
rect 336332 3488 338120 3516
rect 336332 3476 336338 3488
rect 338114 3476 338120 3488
rect 338172 3476 338178 3528
rect 345658 3476 345664 3528
rect 345716 3516 345722 3528
rect 352834 3516 352840 3528
rect 345716 3488 352840 3516
rect 345716 3476 345722 3488
rect 352834 3476 352840 3488
rect 352892 3476 352898 3528
rect 352944 3516 352972 3556
rect 359918 3544 359924 3556
rect 359976 3544 359982 3596
rect 360102 3544 360108 3596
rect 360160 3584 360166 3596
rect 404814 3584 404820 3596
rect 360160 3556 404820 3584
rect 360160 3544 360166 3556
rect 404814 3544 404820 3556
rect 404872 3544 404878 3596
rect 411162 3544 411168 3596
rect 411220 3584 411226 3596
rect 568022 3584 568028 3596
rect 411220 3556 568028 3584
rect 411220 3544 411226 3556
rect 568022 3544 568028 3556
rect 568080 3544 568086 3596
rect 361114 3516 361120 3528
rect 352944 3488 361120 3516
rect 361114 3476 361120 3488
rect 361172 3476 361178 3528
rect 361482 3476 361488 3528
rect 361540 3516 361546 3528
rect 408402 3516 408408 3528
rect 361540 3488 408408 3516
rect 361540 3476 361546 3488
rect 408402 3476 408408 3488
rect 408460 3476 408466 3528
rect 412450 3476 412456 3528
rect 412508 3516 412514 3528
rect 571518 3516 571524 3528
rect 412508 3488 571524 3516
rect 412508 3476 412514 3488
rect 571518 3476 571524 3488
rect 571576 3476 571582 3528
rect 13538 3408 13544 3460
rect 13596 3448 13602 3460
rect 22738 3448 22744 3460
rect 13596 3420 22744 3448
rect 13596 3408 13602 3420
rect 22738 3408 22744 3420
rect 22796 3408 22802 3460
rect 25314 3408 25320 3460
rect 25372 3448 25378 3460
rect 241606 3448 241612 3460
rect 25372 3420 241612 3448
rect 25372 3408 25378 3420
rect 241606 3408 241612 3420
rect 241664 3408 241670 3460
rect 272426 3408 272432 3460
rect 272484 3448 272490 3460
rect 318978 3448 318984 3460
rect 272484 3420 318984 3448
rect 272484 3408 272490 3420
rect 318978 3408 318984 3420
rect 319036 3408 319042 3460
rect 319714 3408 319720 3460
rect 319772 3448 319778 3460
rect 332594 3448 332600 3460
rect 319772 3420 332600 3448
rect 319772 3408 319778 3420
rect 332594 3408 332600 3420
rect 332652 3408 332658 3460
rect 335078 3408 335084 3460
rect 335136 3448 335142 3460
rect 338298 3448 338304 3460
rect 335136 3420 338304 3448
rect 335136 3408 335142 3420
rect 338298 3408 338304 3420
rect 338356 3408 338362 3460
rect 348970 3408 348976 3460
rect 349028 3448 349034 3460
rect 354125 3451 354183 3457
rect 354125 3448 354137 3451
rect 349028 3420 354137 3448
rect 349028 3408 349034 3420
rect 354125 3417 354137 3420
rect 354171 3417 354183 3451
rect 354125 3411 354183 3417
rect 354217 3451 354275 3457
rect 354217 3417 354229 3451
rect 354263 3448 354275 3451
rect 362310 3448 362316 3460
rect 354263 3420 362316 3448
rect 354263 3417 354275 3420
rect 354217 3411 354275 3417
rect 362310 3408 362316 3420
rect 362368 3408 362374 3460
rect 362862 3408 362868 3460
rect 362920 3448 362926 3460
rect 411898 3448 411904 3460
rect 362920 3420 411904 3448
rect 362920 3408 362926 3420
rect 411898 3408 411904 3420
rect 411956 3408 411962 3460
rect 412542 3408 412548 3460
rect 412600 3448 412606 3460
rect 575106 3448 575112 3460
rect 412600 3420 575112 3448
rect 412600 3408 412606 3420
rect 575106 3408 575112 3420
rect 575164 3408 575170 3460
rect 19426 3340 19432 3392
rect 19484 3380 19490 3392
rect 25498 3380 25504 3392
rect 19484 3352 25504 3380
rect 19484 3340 19490 3352
rect 25498 3340 25504 3352
rect 25556 3340 25562 3392
rect 31294 3340 31300 3392
rect 31352 3380 31358 3392
rect 33778 3380 33784 3392
rect 31352 3352 33784 3380
rect 31352 3340 31358 3352
rect 33778 3340 33784 3352
rect 33836 3340 33842 3392
rect 44266 3340 44272 3392
rect 44324 3380 44330 3392
rect 45462 3380 45468 3392
rect 44324 3352 45468 3380
rect 44324 3340 44330 3352
rect 45462 3340 45468 3352
rect 45520 3340 45526 3392
rect 46658 3340 46664 3392
rect 46716 3380 46722 3392
rect 53929 3383 53987 3389
rect 53929 3380 53941 3383
rect 46716 3352 53941 3380
rect 46716 3340 46722 3352
rect 53929 3349 53941 3352
rect 53975 3349 53987 3383
rect 53929 3343 53987 3349
rect 56042 3340 56048 3392
rect 56100 3380 56106 3392
rect 56502 3380 56508 3392
rect 56100 3352 56508 3380
rect 56100 3340 56106 3352
rect 56502 3340 56508 3352
rect 56560 3340 56566 3392
rect 59630 3340 59636 3392
rect 59688 3380 59694 3392
rect 60642 3380 60648 3392
rect 59688 3352 60648 3380
rect 59688 3340 59694 3352
rect 60642 3340 60648 3352
rect 60700 3340 60706 3392
rect 66714 3340 66720 3392
rect 66772 3380 66778 3392
rect 67542 3380 67548 3392
rect 66772 3352 67548 3380
rect 66772 3340 66778 3352
rect 67542 3340 67548 3352
rect 67600 3340 67606 3392
rect 77386 3340 77392 3392
rect 77444 3380 77450 3392
rect 78582 3380 78588 3392
rect 77444 3352 78588 3380
rect 77444 3340 77450 3352
rect 78582 3340 78588 3352
rect 78640 3340 78646 3392
rect 80882 3340 80888 3392
rect 80940 3380 80946 3392
rect 81342 3380 81348 3392
rect 80940 3352 81348 3380
rect 80940 3340 80946 3352
rect 81342 3340 81348 3352
rect 81400 3340 81406 3392
rect 83274 3340 83280 3392
rect 83332 3380 83338 3392
rect 84102 3380 84108 3392
rect 83332 3352 84108 3380
rect 83332 3340 83338 3352
rect 84102 3340 84108 3352
rect 84160 3340 84166 3392
rect 84470 3340 84476 3392
rect 84528 3380 84534 3392
rect 87598 3380 87604 3392
rect 84528 3352 87604 3380
rect 84528 3340 84534 3352
rect 87598 3340 87604 3352
rect 87656 3340 87662 3392
rect 87966 3340 87972 3392
rect 88024 3380 88030 3392
rect 88978 3380 88984 3392
rect 88024 3352 88984 3380
rect 88024 3340 88030 3352
rect 88978 3340 88984 3352
rect 89036 3340 89042 3392
rect 90358 3340 90364 3392
rect 90416 3380 90422 3392
rect 91002 3380 91008 3392
rect 90416 3352 91008 3380
rect 90416 3340 90422 3352
rect 91002 3340 91008 3352
rect 91060 3340 91066 3392
rect 91554 3340 91560 3392
rect 91612 3380 91618 3392
rect 93118 3380 93124 3392
rect 91612 3352 93124 3380
rect 91612 3340 91618 3352
rect 93118 3340 93124 3352
rect 93176 3340 93182 3392
rect 261018 3380 261024 3392
rect 93826 3352 261024 3380
rect 85666 3272 85672 3324
rect 85724 3312 85730 3324
rect 93826 3312 93854 3352
rect 261018 3340 261024 3352
rect 261076 3340 261082 3392
rect 287790 3340 287796 3392
rect 287848 3380 287854 3392
rect 288342 3380 288348 3392
rect 287848 3352 288348 3380
rect 287848 3340 287854 3352
rect 288342 3340 288348 3352
rect 288400 3340 288406 3392
rect 298462 3340 298468 3392
rect 298520 3380 298526 3392
rect 299382 3380 299388 3392
rect 298520 3352 299388 3380
rect 298520 3340 298526 3352
rect 299382 3340 299388 3352
rect 299440 3340 299446 3392
rect 304350 3340 304356 3392
rect 304408 3380 304414 3392
rect 304902 3380 304908 3392
rect 304408 3352 304908 3380
rect 304408 3340 304414 3352
rect 304902 3340 304908 3352
rect 304960 3340 304966 3392
rect 306742 3340 306748 3392
rect 306800 3380 306806 3392
rect 328730 3380 328736 3392
rect 306800 3352 328736 3380
rect 306800 3340 306806 3352
rect 328730 3340 328736 3352
rect 328788 3340 328794 3392
rect 329929 3383 329987 3389
rect 329929 3349 329941 3383
rect 329975 3380 329987 3383
rect 334158 3380 334164 3392
rect 329975 3352 334164 3380
rect 329975 3349 329987 3352
rect 329929 3343 329987 3349
rect 334158 3340 334164 3352
rect 334216 3340 334222 3392
rect 348510 3340 348516 3392
rect 348568 3380 348574 3392
rect 355226 3380 355232 3392
rect 348568 3352 355232 3380
rect 348568 3340 348574 3352
rect 355226 3340 355232 3352
rect 355284 3340 355290 3392
rect 371694 3380 371700 3392
rect 359476 3352 371700 3380
rect 85724 3284 93854 3312
rect 85724 3272 85730 3284
rect 97442 3272 97448 3324
rect 97500 3312 97506 3324
rect 97902 3312 97908 3324
rect 97500 3284 97908 3312
rect 97500 3272 97506 3284
rect 97902 3272 97908 3284
rect 97960 3272 97966 3324
rect 98638 3272 98644 3324
rect 98696 3312 98702 3324
rect 99282 3312 99288 3324
rect 98696 3284 99288 3312
rect 98696 3272 98702 3284
rect 99282 3272 99288 3284
rect 99340 3272 99346 3324
rect 101030 3272 101036 3324
rect 101088 3312 101094 3324
rect 102042 3312 102048 3324
rect 101088 3284 102048 3312
rect 101088 3272 101094 3284
rect 102042 3272 102048 3284
rect 102100 3272 102106 3324
rect 102137 3315 102195 3321
rect 102137 3281 102149 3315
rect 102183 3312 102195 3315
rect 262306 3312 262312 3324
rect 102183 3284 262312 3312
rect 102183 3281 102195 3284
rect 102137 3275 102195 3281
rect 262306 3272 262312 3284
rect 262364 3272 262370 3324
rect 310238 3272 310244 3324
rect 310296 3312 310302 3324
rect 329834 3312 329840 3324
rect 310296 3284 329840 3312
rect 310296 3272 310302 3284
rect 329834 3272 329840 3284
rect 329892 3272 329898 3324
rect 350534 3272 350540 3324
rect 350592 3312 350598 3324
rect 359476 3312 359504 3352
rect 371694 3340 371700 3352
rect 371752 3340 371758 3392
rect 382182 3340 382188 3392
rect 382240 3380 382246 3392
rect 475746 3380 475752 3392
rect 382240 3352 475752 3380
rect 382240 3340 382246 3352
rect 475746 3340 475752 3352
rect 475804 3340 475810 3392
rect 489178 3340 489184 3392
rect 489236 3380 489242 3392
rect 489914 3380 489920 3392
rect 489236 3352 489920 3380
rect 489236 3340 489242 3352
rect 489914 3340 489920 3352
rect 489972 3340 489978 3392
rect 499546 3352 528554 3380
rect 350592 3284 359504 3312
rect 359553 3315 359611 3321
rect 350592 3272 350598 3284
rect 359553 3281 359565 3315
rect 359599 3312 359611 3315
rect 369394 3312 369400 3324
rect 359599 3284 369400 3312
rect 359599 3281 359611 3284
rect 359553 3275 359611 3281
rect 369394 3272 369400 3284
rect 369452 3272 369458 3324
rect 380618 3272 380624 3324
rect 380676 3312 380682 3324
rect 468662 3312 468668 3324
rect 380676 3284 468668 3312
rect 380676 3272 380682 3284
rect 468662 3272 468668 3284
rect 468720 3272 468726 3324
rect 485038 3272 485044 3324
rect 485096 3312 485102 3324
rect 499546 3312 499574 3352
rect 485096 3284 499574 3312
rect 485096 3272 485102 3284
rect 502978 3272 502984 3324
rect 503036 3312 503042 3324
rect 504174 3312 504180 3324
rect 503036 3284 504180 3312
rect 503036 3272 503042 3284
rect 504174 3272 504180 3284
rect 504232 3272 504238 3324
rect 515398 3272 515404 3324
rect 515456 3312 515462 3324
rect 517146 3312 517152 3324
rect 515456 3284 517152 3312
rect 515456 3272 515462 3284
rect 517146 3272 517152 3284
rect 517204 3272 517210 3324
rect 519630 3272 519636 3324
rect 519688 3312 519694 3324
rect 521838 3312 521844 3324
rect 519688 3284 521844 3312
rect 519688 3272 519694 3284
rect 521838 3272 521844 3284
rect 521896 3272 521902 3324
rect 522298 3272 522304 3324
rect 522356 3312 522362 3324
rect 524230 3312 524236 3324
rect 522356 3284 524236 3312
rect 522356 3272 522362 3284
rect 524230 3272 524236 3284
rect 524288 3272 524294 3324
rect 528526 3312 528554 3352
rect 530578 3340 530584 3392
rect 530636 3380 530642 3392
rect 531314 3380 531320 3392
rect 530636 3352 531320 3380
rect 530636 3340 530642 3352
rect 531314 3340 531320 3352
rect 531372 3340 531378 3392
rect 533338 3340 533344 3392
rect 533396 3380 533402 3392
rect 534902 3380 534908 3392
rect 533396 3352 534908 3380
rect 533396 3340 533402 3352
rect 534902 3340 534908 3352
rect 534960 3340 534966 3392
rect 534997 3383 535055 3389
rect 534997 3349 535009 3383
rect 535043 3380 535055 3383
rect 539594 3380 539600 3392
rect 535043 3352 539600 3380
rect 535043 3349 535055 3352
rect 534997 3343 535055 3349
rect 539594 3340 539600 3352
rect 539652 3340 539658 3392
rect 540238 3340 540244 3392
rect 540296 3380 540302 3392
rect 541986 3380 541992 3392
rect 540296 3352 541992 3380
rect 540296 3340 540302 3352
rect 541986 3340 541992 3352
rect 542044 3340 542050 3392
rect 532510 3312 532516 3324
rect 528526 3284 532516 3312
rect 532510 3272 532516 3284
rect 532568 3272 532574 3324
rect 92750 3204 92756 3256
rect 92808 3244 92814 3256
rect 262490 3244 262496 3256
rect 92808 3216 262496 3244
rect 92808 3204 92814 3216
rect 262490 3204 262496 3216
rect 262548 3204 262554 3256
rect 311434 3204 311440 3256
rect 311492 3244 311498 3256
rect 329926 3244 329932 3256
rect 311492 3216 329932 3244
rect 311492 3204 311498 3216
rect 329926 3204 329932 3216
rect 329984 3204 329990 3256
rect 331490 3244 331496 3256
rect 330036 3216 331496 3244
rect 57238 3136 57244 3188
rect 57296 3176 57302 3188
rect 61378 3176 61384 3188
rect 57296 3148 61384 3176
rect 57296 3136 57302 3148
rect 61378 3136 61384 3148
rect 61436 3136 61442 3188
rect 93946 3136 93952 3188
rect 94004 3176 94010 3188
rect 95050 3176 95056 3188
rect 94004 3148 95056 3176
rect 94004 3136 94010 3148
rect 95050 3136 95056 3148
rect 95108 3136 95114 3188
rect 96246 3136 96252 3188
rect 96304 3176 96310 3188
rect 263778 3176 263784 3188
rect 96304 3148 263784 3176
rect 96304 3136 96310 3148
rect 263778 3136 263784 3148
rect 263836 3136 263842 3188
rect 312630 3136 312636 3188
rect 312688 3176 312694 3188
rect 330036 3176 330064 3216
rect 331490 3204 331496 3216
rect 331548 3204 331554 3256
rect 349062 3204 349068 3256
rect 349120 3244 349126 3256
rect 365806 3244 365812 3256
rect 349120 3216 365812 3244
rect 349120 3204 349126 3216
rect 365806 3204 365812 3216
rect 365864 3204 365870 3256
rect 377766 3204 377772 3256
rect 377824 3244 377830 3256
rect 461578 3244 461584 3256
rect 377824 3216 461584 3244
rect 377824 3204 377830 3216
rect 461578 3204 461584 3216
rect 461636 3204 461642 3256
rect 526438 3204 526444 3256
rect 526496 3244 526502 3256
rect 527818 3244 527824 3256
rect 526496 3216 527824 3244
rect 526496 3204 526502 3216
rect 527818 3204 527824 3216
rect 527876 3204 527882 3256
rect 312688 3148 330064 3176
rect 312688 3136 312694 3148
rect 330386 3136 330392 3188
rect 330444 3176 330450 3188
rect 333238 3176 333244 3188
rect 330444 3148 333244 3176
rect 330444 3136 330450 3148
rect 333238 3136 333244 3148
rect 333296 3136 333302 3188
rect 342162 3136 342168 3188
rect 342220 3176 342226 3188
rect 344554 3176 344560 3188
rect 342220 3148 344560 3176
rect 342220 3136 342226 3148
rect 344554 3136 344560 3148
rect 344612 3136 344618 3188
rect 347038 3136 347044 3188
rect 347096 3176 347102 3188
rect 354030 3176 354036 3188
rect 347096 3148 354036 3176
rect 347096 3136 347102 3148
rect 354030 3136 354036 3148
rect 354088 3136 354094 3188
rect 354125 3179 354183 3185
rect 354125 3145 354137 3179
rect 354171 3176 354183 3179
rect 359553 3179 359611 3185
rect 359553 3176 359565 3179
rect 354171 3148 359565 3176
rect 354171 3145 354183 3148
rect 354125 3139 354183 3145
rect 359553 3145 359565 3148
rect 359599 3145 359611 3179
rect 364610 3176 364616 3188
rect 359553 3139 359611 3145
rect 364306 3148 364616 3176
rect 89162 3068 89168 3120
rect 89220 3108 89226 3120
rect 102137 3111 102195 3117
rect 102137 3108 102149 3111
rect 89220 3080 102149 3108
rect 89220 3068 89226 3080
rect 102137 3077 102149 3080
rect 102183 3077 102195 3111
rect 102137 3071 102195 3077
rect 102226 3068 102232 3120
rect 102284 3108 102290 3120
rect 104158 3108 104164 3120
rect 102284 3080 104164 3108
rect 102284 3068 102290 3080
rect 104158 3068 104164 3080
rect 104216 3068 104222 3120
rect 105722 3068 105728 3120
rect 105780 3108 105786 3120
rect 106182 3108 106188 3120
rect 105780 3080 106188 3108
rect 105780 3068 105786 3080
rect 106182 3068 106188 3080
rect 106240 3068 106246 3120
rect 106918 3068 106924 3120
rect 106976 3108 106982 3120
rect 107562 3108 107568 3120
rect 106976 3080 107568 3108
rect 106976 3068 106982 3080
rect 107562 3068 107568 3080
rect 107620 3068 107626 3120
rect 108114 3068 108120 3120
rect 108172 3108 108178 3120
rect 108942 3108 108948 3120
rect 108172 3080 108948 3108
rect 108172 3068 108178 3080
rect 108942 3068 108948 3080
rect 109000 3068 109006 3120
rect 109310 3068 109316 3120
rect 109368 3108 109374 3120
rect 111058 3108 111064 3120
rect 109368 3080 111064 3108
rect 109368 3068 109374 3080
rect 111058 3068 111064 3080
rect 111116 3068 111122 3120
rect 111153 3111 111211 3117
rect 111153 3077 111165 3111
rect 111199 3108 111211 3111
rect 265250 3108 265256 3120
rect 111199 3080 265256 3108
rect 111199 3077 111211 3080
rect 111153 3071 111211 3077
rect 265250 3068 265256 3080
rect 265308 3068 265314 3120
rect 313826 3068 313832 3120
rect 313884 3108 313890 3120
rect 331398 3108 331404 3120
rect 313884 3080 331404 3108
rect 313884 3068 313890 3080
rect 331398 3068 331404 3080
rect 331456 3068 331462 3120
rect 338666 3068 338672 3120
rect 338724 3108 338730 3120
rect 339586 3108 339592 3120
rect 338724 3080 339592 3108
rect 338724 3068 338730 3080
rect 339586 3068 339592 3080
rect 339644 3068 339650 3120
rect 349798 3068 349804 3120
rect 349856 3108 349862 3120
rect 357526 3108 357532 3120
rect 349856 3080 357532 3108
rect 349856 3068 349862 3080
rect 357526 3068 357532 3080
rect 357584 3068 357590 3120
rect 27706 3000 27712 3052
rect 27764 3040 27770 3052
rect 29638 3040 29644 3052
rect 27764 3012 29644 3040
rect 27764 3000 27770 3012
rect 29638 3000 29644 3012
rect 29696 3000 29702 3052
rect 73798 3000 73804 3052
rect 73856 3040 73862 3052
rect 74442 3040 74448 3052
rect 73856 3012 74448 3040
rect 73856 3000 73862 3012
rect 74442 3000 74448 3012
rect 74500 3000 74506 3052
rect 103330 3000 103336 3052
rect 103388 3040 103394 3052
rect 266630 3040 266636 3052
rect 103388 3012 266636 3040
rect 103388 3000 103394 3012
rect 266630 3000 266636 3012
rect 266688 3000 266694 3052
rect 296070 3000 296076 3052
rect 296128 3040 296134 3052
rect 296622 3040 296628 3052
rect 296128 3012 296628 3040
rect 296128 3000 296134 3012
rect 296622 3000 296628 3012
rect 296680 3000 296686 3052
rect 315022 3000 315028 3052
rect 315080 3040 315086 3052
rect 331214 3040 331220 3052
rect 315080 3012 331220 3040
rect 315080 3000 315086 3012
rect 331214 3000 331220 3012
rect 331272 3000 331278 3052
rect 337470 3000 337476 3052
rect 337528 3040 337534 3052
rect 338206 3040 338212 3052
rect 337528 3012 338212 3040
rect 337528 3000 337534 3012
rect 338206 3000 338212 3012
rect 338264 3000 338270 3052
rect 348418 3000 348424 3052
rect 348476 3040 348482 3052
rect 364306 3040 364334 3148
rect 364610 3136 364616 3148
rect 364668 3136 364674 3188
rect 375098 3136 375104 3188
rect 375156 3176 375162 3188
rect 454494 3176 454500 3188
rect 375156 3148 454500 3176
rect 375156 3136 375162 3148
rect 454494 3136 454500 3148
rect 454552 3136 454558 3188
rect 456794 3136 456800 3188
rect 456852 3176 456858 3188
rect 458082 3176 458088 3188
rect 456852 3148 458088 3176
rect 456852 3136 456858 3148
rect 458082 3136 458088 3148
rect 458140 3136 458146 3188
rect 512638 3136 512644 3188
rect 512696 3176 512702 3188
rect 513558 3176 513564 3188
rect 512696 3148 513564 3176
rect 512696 3136 512702 3148
rect 513558 3136 513564 3148
rect 513616 3136 513622 3188
rect 373902 3068 373908 3120
rect 373960 3108 373966 3120
rect 447410 3108 447416 3120
rect 373960 3080 447416 3108
rect 373960 3068 373966 3080
rect 447410 3068 447416 3080
rect 447468 3068 447474 3120
rect 348476 3012 364334 3040
rect 348476 3000 348482 3012
rect 371142 3000 371148 3052
rect 371200 3040 371206 3052
rect 440326 3040 440332 3052
rect 371200 3012 440332 3040
rect 371200 3000 371206 3012
rect 440326 3000 440332 3012
rect 440384 3000 440390 3052
rect 99834 2932 99840 2984
rect 99892 2972 99898 2984
rect 99892 2944 103514 2972
rect 99892 2932 99898 2944
rect 9950 2864 9956 2916
rect 10008 2904 10014 2916
rect 14458 2904 14464 2916
rect 10008 2876 14464 2904
rect 10008 2864 10014 2876
rect 14458 2864 14464 2876
rect 14516 2864 14522 2916
rect 103486 2904 103514 2944
rect 110506 2932 110512 2984
rect 110564 2972 110570 2984
rect 267918 2972 267924 2984
rect 110564 2944 267924 2972
rect 110564 2932 110570 2944
rect 267918 2932 267924 2944
rect 267976 2932 267982 2984
rect 317322 2932 317328 2984
rect 317380 2972 317386 2984
rect 332778 2972 332784 2984
rect 317380 2944 332784 2972
rect 317380 2932 317386 2944
rect 332778 2932 332784 2944
rect 332836 2932 332842 2984
rect 355962 2932 355968 2984
rect 356020 2972 356026 2984
rect 363785 2975 363843 2981
rect 363785 2972 363797 2975
rect 356020 2944 363797 2972
rect 356020 2932 356026 2944
rect 363785 2941 363797 2944
rect 363831 2941 363843 2975
rect 363785 2935 363843 2941
rect 369762 2932 369768 2984
rect 369820 2972 369826 2984
rect 433242 2972 433248 2984
rect 369820 2944 433248 2972
rect 369820 2932 369826 2944
rect 433242 2932 433248 2944
rect 433300 2932 433306 2984
rect 111153 2907 111211 2913
rect 111153 2904 111165 2907
rect 103486 2876 111165 2904
rect 111153 2873 111165 2876
rect 111199 2873 111211 2907
rect 111153 2867 111211 2873
rect 114002 2864 114008 2916
rect 114060 2904 114066 2916
rect 114462 2904 114468 2916
rect 114060 2876 114468 2904
rect 114060 2864 114066 2876
rect 114462 2864 114468 2876
rect 114520 2864 114526 2916
rect 115198 2864 115204 2916
rect 115256 2904 115262 2916
rect 115842 2904 115848 2916
rect 115256 2876 115848 2904
rect 115256 2864 115262 2876
rect 115842 2864 115848 2876
rect 115900 2864 115906 2916
rect 116394 2864 116400 2916
rect 116452 2904 116458 2916
rect 117222 2904 117228 2916
rect 116452 2876 117228 2904
rect 116452 2864 116458 2876
rect 117222 2864 117228 2876
rect 117280 2864 117286 2916
rect 118786 2864 118792 2916
rect 118844 2904 118850 2916
rect 119798 2904 119804 2916
rect 118844 2876 119804 2904
rect 118844 2864 118850 2876
rect 119798 2864 119804 2876
rect 119856 2864 119862 2916
rect 270770 2904 270776 2916
rect 120092 2876 270776 2904
rect 117590 2796 117596 2848
rect 117648 2836 117654 2848
rect 120092 2836 120120 2876
rect 270770 2864 270776 2876
rect 270828 2864 270834 2916
rect 276014 2864 276020 2916
rect 276072 2904 276078 2916
rect 277302 2904 277308 2916
rect 276072 2876 277308 2904
rect 276072 2864 276078 2876
rect 277302 2864 277308 2876
rect 277360 2864 277366 2916
rect 318518 2864 318524 2916
rect 318576 2904 318582 2916
rect 332870 2904 332876 2916
rect 318576 2876 332876 2904
rect 318576 2864 318582 2876
rect 332870 2864 332876 2876
rect 332928 2864 332934 2916
rect 365622 2864 365628 2916
rect 365680 2904 365686 2916
rect 422570 2904 422576 2916
rect 365680 2876 422576 2904
rect 365680 2864 365686 2876
rect 422570 2864 422576 2876
rect 422628 2864 422634 2916
rect 117648 2808 120120 2836
rect 117648 2796 117654 2808
rect 121086 2796 121092 2848
rect 121144 2836 121150 2848
rect 272058 2836 272064 2848
rect 121144 2808 272064 2836
rect 121144 2796 121150 2808
rect 272058 2796 272064 2808
rect 272116 2796 272122 2848
rect 316218 2796 316224 2848
rect 316276 2836 316282 2848
rect 331306 2836 331312 2848
rect 316276 2808 331312 2836
rect 316276 2796 316282 2808
rect 331306 2796 331312 2808
rect 331364 2796 331370 2848
rect 364242 2796 364248 2848
rect 364300 2836 364306 2848
rect 415486 2836 415492 2848
rect 364300 2808 415492 2836
rect 364300 2796 364306 2808
rect 415486 2796 415492 2808
rect 415544 2796 415550 2848
<< via1 >>
rect 317328 700952 317380 701004
rect 429844 700952 429896 701004
rect 202788 700884 202840 700936
rect 331312 700884 331364 700936
rect 313188 700816 313240 700868
rect 462320 700816 462372 700868
rect 315948 700748 316000 700800
rect 478512 700748 478564 700800
rect 311808 700680 311860 700732
rect 494796 700680 494848 700732
rect 137836 700612 137888 700664
rect 336740 700612 336792 700664
rect 309048 700544 309100 700596
rect 527180 700544 527232 700596
rect 105452 700476 105504 700528
rect 106188 700476 106240 700528
rect 310428 700476 310480 700528
rect 543464 700476 543516 700528
rect 40500 700408 40552 700460
rect 41328 700408 41380 700460
rect 307668 700408 307720 700460
rect 559656 700408 559708 700460
rect 72976 700340 73028 700392
rect 340880 700340 340932 700392
rect 8116 700272 8168 700324
rect 345020 700272 345072 700324
rect 320088 700204 320140 700256
rect 413652 700204 413704 700256
rect 318708 700136 318760 700188
rect 397460 700136 397512 700188
rect 267648 700068 267700 700120
rect 327080 700068 327132 700120
rect 321468 700000 321520 700052
rect 364984 700000 365036 700052
rect 324228 699932 324280 699984
rect 348792 699932 348844 699984
rect 322848 699864 322900 699916
rect 332508 699864 332560 699916
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 170312 699660 170364 699712
rect 171048 699660 171100 699712
rect 235172 699660 235224 699712
rect 235908 699660 235960 699712
rect 300124 699660 300176 699712
rect 300768 699660 300820 699712
rect 304908 696940 304960 696992
rect 580172 696940 580224 696992
rect 306288 683136 306340 683188
rect 580172 683136 580224 683188
rect 302148 670692 302200 670744
rect 580172 670692 580224 670744
rect 3148 656888 3200 656940
rect 350540 656888 350592 656940
rect 299388 643084 299440 643136
rect 580172 643084 580224 643136
rect 300676 630640 300728 630692
rect 580172 630640 580224 630692
rect 2964 618264 3016 618316
rect 333244 618264 333296 618316
rect 298008 616836 298060 616888
rect 580172 616836 580224 616888
rect 3332 605820 3384 605872
rect 354680 605820 354732 605872
rect 295248 590656 295300 590708
rect 579804 590656 579856 590708
rect 296628 576852 296680 576904
rect 580172 576852 580224 576904
rect 3332 565836 3384 565888
rect 338764 565836 338816 565888
rect 293868 563048 293920 563100
rect 579804 563048 579856 563100
rect 3332 553392 3384 553444
rect 360200 553392 360252 553444
rect 289728 536800 289780 536852
rect 580172 536800 580224 536852
rect 291108 524424 291160 524476
rect 580172 524424 580224 524476
rect 3332 514768 3384 514820
rect 342904 514768 342956 514820
rect 288348 510620 288400 510672
rect 580172 510620 580224 510672
rect 3240 500964 3292 501016
rect 364340 500964 364392 501016
rect 285588 484372 285640 484424
rect 580172 484372 580224 484424
rect 286968 470568 287020 470620
rect 579988 470568 580040 470620
rect 3516 462340 3568 462392
rect 348516 462340 348568 462392
rect 154488 460844 154540 460896
rect 338120 460844 338172 460896
rect 338764 460844 338816 460896
rect 361764 460844 361816 460896
rect 106188 460776 106240 460828
rect 339684 460776 339736 460828
rect 89628 460708 89680 460760
rect 342812 460708 342864 460760
rect 342904 460708 342956 460760
rect 366456 460708 366508 460760
rect 41328 460640 41380 460692
rect 344376 460640 344428 460692
rect 24768 460572 24820 460624
rect 347780 460572 347832 460624
rect 348516 460572 348568 460624
rect 371240 460572 371292 460624
rect 3424 460504 3476 460556
rect 349160 460504 349212 460556
rect 3608 460436 3660 460488
rect 352288 460436 352340 460488
rect 3700 460368 3752 460420
rect 353852 460368 353904 460420
rect 3792 460300 3844 460352
rect 358820 460300 358872 460352
rect 3884 460232 3936 460284
rect 363328 460232 363380 460284
rect 3976 460164 4028 460216
rect 368112 460164 368164 460216
rect 171048 460096 171100 460148
rect 334900 460096 334952 460148
rect 219348 460028 219400 460080
rect 235908 459960 235960 460012
rect 330208 459960 330260 460012
rect 333244 460028 333296 460080
rect 356980 460028 357032 460080
rect 333336 459960 333388 460012
rect 284208 459892 284260 459944
rect 328552 459892 328604 459944
rect 300768 459756 300820 459808
rect 325700 459824 325752 459876
rect 281448 459688 281500 459740
rect 285036 459620 285088 459672
rect 285588 459620 285640 459672
rect 292948 459688 293000 459740
rect 293868 459688 293920 459740
rect 294512 459688 294564 459740
rect 295248 459688 295300 459740
rect 296076 459688 296128 459740
rect 296628 459688 296680 459740
rect 303988 459688 304040 459740
rect 304908 459688 304960 459740
rect 305552 459688 305604 459740
rect 306288 459688 306340 459740
rect 307116 459688 307168 459740
rect 307668 459688 307720 459740
rect 315028 459688 315080 459740
rect 315948 459688 316000 459740
rect 316592 459688 316644 459740
rect 317328 459688 317380 459740
rect 318156 459688 318208 459740
rect 318708 459688 318760 459740
rect 556804 459620 556856 459672
rect 272340 459552 272392 459604
rect 555424 459552 555476 459604
rect 255044 458804 255096 458856
rect 580264 458804 580316 458856
rect 278688 458668 278740 458720
rect 418804 458668 418856 458720
rect 280068 458600 280120 458652
rect 428464 458600 428516 458652
rect 228364 458532 228416 458584
rect 379152 458532 379204 458584
rect 270408 458464 270460 458516
rect 421656 458464 421708 458516
rect 222844 458396 222896 458448
rect 375932 458396 375984 458448
rect 277032 458328 277084 458380
rect 429844 458328 429896 458380
rect 232596 458260 232648 458312
rect 391940 458260 391992 458312
rect 3424 458192 3476 458244
rect 373126 458192 373178 458244
rect 233884 457376 233936 457428
rect 239220 457419 239272 457428
rect 239220 457385 239229 457419
rect 239229 457385 239263 457419
rect 239263 457385 239272 457419
rect 239220 457376 239272 457385
rect 273996 457419 274048 457428
rect 273996 457385 274005 457419
rect 274005 457385 274039 457419
rect 274039 457385 274048 457419
rect 273996 457376 274048 457385
rect 275560 457419 275612 457428
rect 275560 457385 275569 457419
rect 275569 457385 275603 457419
rect 275603 457385 275612 457419
rect 275560 457376 275612 457385
rect 283472 457419 283524 457428
rect 283472 457385 283481 457419
rect 283481 457385 283515 457419
rect 283515 457385 283524 457419
rect 283472 457376 283524 457385
rect 369860 457308 369912 457360
rect 231124 457240 231176 457292
rect 374368 457308 374420 457360
rect 377588 457351 377640 457360
rect 377588 457317 377597 457351
rect 377597 457317 377631 457351
rect 377631 457317 377640 457351
rect 377588 457308 377640 457317
rect 380900 457351 380952 457360
rect 380900 457317 380909 457351
rect 380909 457317 380943 457351
rect 380943 457317 380952 457351
rect 380900 457308 380952 457317
rect 407580 457351 407632 457360
rect 407580 457317 407589 457351
rect 407589 457317 407623 457351
rect 407623 457317 407632 457351
rect 407580 457308 407632 457317
rect 417424 457172 417476 457224
rect 425704 457104 425756 457156
rect 224224 457036 224276 457088
rect 226984 456968 227036 457020
rect 431224 456900 431276 456952
rect 579804 456832 579856 456884
rect 4804 456764 4856 456816
rect 3332 449828 3384 449880
rect 233884 449828 233936 449880
rect 428464 431876 428516 431928
rect 580172 431876 580224 431928
rect 556804 419432 556856 419484
rect 580172 419432 580224 419484
rect 3424 411204 3476 411256
rect 222844 411204 222896 411256
rect 418804 405628 418856 405680
rect 579620 405628 579672 405680
rect 3240 398760 3292 398812
rect 231124 398760 231176 398812
rect 425704 379448 425756 379500
rect 580172 379448 580224 379500
rect 2780 371424 2832 371476
rect 4804 371424 4856 371476
rect 429844 365644 429896 365696
rect 580172 365644 580224 365696
rect 3332 358708 3384 358760
rect 224224 358708 224276 358760
rect 417424 353200 417476 353252
rect 580172 353200 580224 353252
rect 3148 346332 3200 346384
rect 228364 346332 228416 346384
rect 220084 336676 220136 336728
rect 288440 336676 288492 336728
rect 289820 336676 289872 336728
rect 291568 336676 291620 336728
rect 292948 336676 293000 336728
rect 300492 336676 300544 336728
rect 301320 336676 301372 336728
rect 304908 336676 304960 336728
rect 328552 336676 328604 336728
rect 339500 336676 339552 336728
rect 339776 336676 339828 336728
rect 342720 336676 342772 336728
rect 343456 336676 343508 336728
rect 343548 336676 343600 336728
rect 344284 336676 344336 336728
rect 347044 336676 347096 336728
rect 347596 336676 347648 336728
rect 354036 336676 354088 336728
rect 354496 336676 354548 336728
rect 355048 336676 355100 336728
rect 355784 336676 355836 336728
rect 356520 336676 356572 336728
rect 357164 336676 357216 336728
rect 357992 336676 358044 336728
rect 358728 336676 358780 336728
rect 359464 336676 359516 336728
rect 359924 336676 359976 336728
rect 360936 336676 360988 336728
rect 361396 336676 361448 336728
rect 362592 336676 362644 336728
rect 362868 336676 362920 336728
rect 363512 336676 363564 336728
rect 364248 336676 364300 336728
rect 370412 336676 370464 336728
rect 435364 336676 435416 336728
rect 215944 336608 215996 336660
rect 292212 336608 292264 336660
rect 292488 336608 292540 336660
rect 295432 336608 295484 336660
rect 296536 336608 296588 336660
rect 296904 336608 296956 336660
rect 300768 336608 300820 336660
rect 327540 336608 327592 336660
rect 341248 336608 341300 336660
rect 342444 336608 342496 336660
rect 349620 336608 349672 336660
rect 353944 336608 353996 336660
rect 355692 336608 355744 336660
rect 355968 336608 356020 336660
rect 359096 336608 359148 336660
rect 360016 336608 360068 336660
rect 362040 336608 362092 336660
rect 362684 336608 362736 336660
rect 369768 336608 369820 336660
rect 436100 336608 436152 336660
rect 214564 336540 214616 336592
rect 293316 336540 293368 336592
rect 296628 336540 296680 336592
rect 326160 336540 326212 336592
rect 345572 336540 345624 336592
rect 349804 336540 349856 336592
rect 372252 336540 372304 336592
rect 443000 336540 443052 336592
rect 209044 336472 209096 336524
rect 296720 336472 296772 336524
rect 299388 336472 299440 336524
rect 327080 336472 327132 336524
rect 329104 336472 329156 336524
rect 333980 336472 334032 336524
rect 348516 336472 348568 336524
rect 363604 336472 363656 336524
rect 373356 336472 373408 336524
rect 373908 336472 373960 336524
rect 374828 336472 374880 336524
rect 375196 336472 375248 336524
rect 375932 336472 375984 336524
rect 376668 336472 376720 336524
rect 377036 336472 377088 336524
rect 377864 336472 377916 336524
rect 380256 336472 380308 336524
rect 380716 336472 380768 336524
rect 382004 336472 382056 336524
rect 382188 336472 382240 336524
rect 449900 336472 449952 336524
rect 125508 336404 125560 336456
rect 114468 336336 114520 336388
rect 269948 336336 270000 336388
rect 271788 336404 271840 336456
rect 272800 336404 272852 336456
rect 276020 336404 276072 336456
rect 277860 336404 277912 336456
rect 279792 336404 279844 336456
rect 282644 336404 282696 336456
rect 283380 336404 283432 336456
rect 294420 336404 294472 336456
rect 323584 336404 323636 336456
rect 347412 336404 347464 336456
rect 367836 336404 367888 336456
rect 379888 336404 379940 336456
rect 380624 336404 380676 336456
rect 456800 336404 456852 336456
rect 273260 336336 273312 336388
rect 277308 336336 277360 336388
rect 319904 336336 319956 336388
rect 347688 336336 347740 336388
rect 348424 336336 348476 336388
rect 354404 336336 354456 336388
rect 370504 336336 370556 336388
rect 374460 336336 374512 336388
rect 378876 336336 378928 336388
rect 465080 336336 465132 336388
rect 107568 336268 107620 336320
rect 267832 336268 267884 336320
rect 279056 336268 279108 336320
rect 282184 336268 282236 336320
rect 283104 336268 283156 336320
rect 321560 336268 321612 336320
rect 348884 336268 348936 336320
rect 367376 336268 367428 336320
rect 368204 336268 368256 336320
rect 57244 336200 57296 336252
rect 251272 336200 251324 336252
rect 259460 336200 259512 336252
rect 261484 336200 261536 336252
rect 264888 336200 264940 336252
rect 265164 336200 265216 336252
rect 269120 336200 269172 336252
rect 271880 336200 271932 336252
rect 274548 336200 274600 336252
rect 319260 336200 319312 336252
rect 327724 336200 327776 336252
rect 328460 336200 328512 336252
rect 341616 336200 341668 336252
rect 342168 336200 342220 336252
rect 346676 336200 346728 336252
rect 347688 336200 347740 336252
rect 352196 336200 352248 336252
rect 371792 336200 371844 336252
rect 373724 336200 373776 336252
rect 374276 336200 374328 336252
rect 51724 336132 51776 336184
rect 247960 336132 248012 336184
rect 267648 336132 267700 336184
rect 317052 336132 317104 336184
rect 351460 336132 351512 336184
rect 50344 336064 50396 336116
rect 245844 336064 245896 336116
rect 270408 336064 270460 336116
rect 318156 336064 318208 336116
rect 344100 336064 344152 336116
rect 345664 336064 345716 336116
rect 348148 336064 348200 336116
rect 349068 336064 349120 336116
rect 351092 336064 351144 336116
rect 351828 336064 351880 336116
rect 352564 336064 352616 336116
rect 353208 336064 353260 336116
rect 358084 336132 358136 336184
rect 363880 336132 363932 336184
rect 375472 336064 375524 336116
rect 376576 336200 376628 336252
rect 381728 336268 381780 336320
rect 468484 336268 468536 336320
rect 380808 336200 380860 336252
rect 471980 336200 472032 336252
rect 383476 336132 383528 336184
rect 475384 336132 475436 336184
rect 382924 336064 382976 336116
rect 383200 336064 383252 336116
rect 478880 336064 478932 336116
rect 35164 335996 35216 336048
rect 243636 335996 243688 336048
rect 263508 335996 263560 336048
rect 316040 335996 316092 336048
rect 316684 335996 316736 336048
rect 327264 335996 327316 336048
rect 328368 335996 328420 336048
rect 336004 335996 336056 336048
rect 344836 335996 344888 336048
rect 348516 335996 348568 336048
rect 353668 335996 353720 336048
rect 382464 335996 382516 336048
rect 383936 335996 383988 336048
rect 384856 335996 384908 336048
rect 387248 335996 387300 336048
rect 387708 335996 387760 336048
rect 388352 335996 388404 336048
rect 389088 335996 389140 336048
rect 389456 335996 389508 336048
rect 390192 335996 390244 336048
rect 392676 335996 392728 336048
rect 393136 335996 393188 336048
rect 395344 335996 395396 336048
rect 397828 335996 397880 336048
rect 398564 335996 398616 336048
rect 402244 335996 402296 336048
rect 402704 335996 402756 336048
rect 497464 335996 497516 336048
rect 204904 335928 204956 335980
rect 276848 335928 276900 335980
rect 281356 335928 281408 335980
rect 286416 335928 286468 335980
rect 315212 335928 315264 335980
rect 346308 335928 346360 335980
rect 347136 335928 347188 335980
rect 356888 335928 356940 335980
rect 357348 335928 357400 335980
rect 369308 335928 369360 335980
rect 432604 335928 432656 335980
rect 224224 335860 224276 335912
rect 291200 335860 291252 335912
rect 291936 335860 291988 335912
rect 311900 335860 311952 335912
rect 333244 335860 333296 335912
rect 336740 335860 336792 335912
rect 364616 335860 364668 335912
rect 372988 335860 373040 335912
rect 374644 335860 374696 335912
rect 429200 335860 429252 335912
rect 233884 335792 233936 335844
rect 300216 335792 300268 335844
rect 336004 335792 336056 335844
rect 337476 335792 337528 335844
rect 361028 335792 361080 335844
rect 361488 335792 361540 335844
rect 366456 335792 366508 335844
rect 367008 335792 367060 335844
rect 367468 335792 367520 335844
rect 368296 335792 368348 335844
rect 428464 335792 428516 335844
rect 222844 335724 222896 335776
rect 287796 335724 287848 335776
rect 289084 335724 289136 335776
rect 313004 335724 313056 335776
rect 366824 335724 366876 335776
rect 425060 335724 425112 335776
rect 213184 335656 213236 335708
rect 273904 335656 273956 335708
rect 288348 335656 288400 335708
rect 295984 335656 296036 335708
rect 228364 335588 228416 335640
rect 288900 335588 288952 335640
rect 296444 335588 296496 335640
rect 298100 335588 298152 335640
rect 310520 335656 310572 335708
rect 310796 335656 310848 335708
rect 360568 335656 360620 335708
rect 361304 335656 361356 335708
rect 368940 335656 368992 335708
rect 369768 335656 369820 335708
rect 314936 335588 314988 335640
rect 366088 335588 366140 335640
rect 413192 335656 413244 335708
rect 413836 335656 413888 335708
rect 414756 335656 414808 335708
rect 415308 335656 415360 335708
rect 231124 335520 231176 335572
rect 285680 335520 285732 335572
rect 344468 335520 344520 335572
rect 346952 335520 347004 335572
rect 352932 335520 352984 335572
rect 353116 335520 353168 335572
rect 364984 335520 365036 335572
rect 371884 335520 371936 335572
rect 372344 335520 372396 335572
rect 414664 335588 414716 335640
rect 415216 335588 415268 335640
rect 417516 335520 417568 335572
rect 232504 335452 232556 335504
rect 282368 335452 282420 335504
rect 366916 335452 366968 335504
rect 418804 335452 418856 335504
rect 233976 335384 234028 335436
rect 273536 335384 273588 335436
rect 341984 335384 342036 335436
rect 345204 335384 345256 335436
rect 350080 335384 350132 335436
rect 350356 335384 350408 335436
rect 357440 335384 357492 335436
rect 401876 335384 401928 335436
rect 402612 335384 402664 335436
rect 403992 335384 404044 335436
rect 404268 335384 404320 335436
rect 404728 335384 404780 335436
rect 405280 335384 405332 335436
rect 405372 335384 405424 335436
rect 405556 335384 405608 335436
rect 406568 335384 406620 335436
rect 406844 335384 406896 335436
rect 407672 335384 407724 335436
rect 408316 335384 408368 335436
rect 409512 335384 409564 335436
rect 409788 335384 409840 335436
rect 410708 335384 410760 335436
rect 411076 335384 411128 335436
rect 412088 335384 412140 335436
rect 412364 335384 412416 335436
rect 418160 335384 418212 335436
rect 274456 335316 274508 335368
rect 278780 335316 278832 335368
rect 179328 335248 179380 335300
rect 290004 335316 290056 335368
rect 332508 335316 332560 335368
rect 337108 335316 337160 335368
rect 344928 335316 344980 335368
rect 345756 335316 345808 335368
rect 355416 335316 355468 335368
rect 388444 335316 388496 335368
rect 388812 335316 388864 335368
rect 403256 335316 403308 335368
rect 404176 335316 404228 335368
rect 405096 335316 405148 335368
rect 405648 335316 405700 335368
rect 406200 335316 406252 335368
rect 407028 335316 407080 335368
rect 408776 335316 408828 335368
rect 409604 335316 409656 335368
rect 410248 335316 410300 335368
rect 410984 335316 411036 335368
rect 411720 335316 411772 335368
rect 412456 335316 412508 335368
rect 421564 335316 421616 335368
rect 388996 335248 389048 335300
rect 483020 335248 483072 335300
rect 169668 335180 169720 335232
rect 286692 335180 286744 335232
rect 384304 335180 384356 335232
rect 481640 335180 481692 335232
rect 161388 335112 161440 335164
rect 284484 335112 284536 335164
rect 391940 335112 391992 335164
rect 490012 335112 490064 335164
rect 144828 335044 144880 335096
rect 276020 335044 276072 335096
rect 390100 335044 390152 335096
rect 500960 335044 501012 335096
rect 147588 334976 147640 335028
rect 280252 334976 280304 335028
rect 392308 334976 392360 335028
rect 507860 334976 507912 335028
rect 140688 334908 140740 334960
rect 277952 334908 278004 334960
rect 393780 334908 393832 334960
rect 512644 334908 512696 334960
rect 86868 334840 86920 334892
rect 259460 334840 259512 334892
rect 395896 334840 395948 334892
rect 520280 334840 520332 334892
rect 87604 334772 87656 334824
rect 260932 334772 260984 334824
rect 398196 334772 398248 334824
rect 526444 334772 526496 334824
rect 54484 334704 54536 334756
rect 247592 334704 247644 334756
rect 397092 334704 397144 334756
rect 522304 334704 522356 334756
rect 29644 334636 29696 334688
rect 243268 334636 243320 334688
rect 398472 334636 398524 334688
rect 528560 334636 528612 334688
rect 22744 334568 22796 334620
rect 238852 334568 238904 334620
rect 402520 334568 402572 334620
rect 540244 334568 540296 334620
rect 197268 334500 197320 334552
rect 292488 334500 292540 334552
rect 374276 334500 374328 334552
rect 448520 334500 448572 334552
rect 202788 334432 202840 334484
rect 296536 334432 296588 334484
rect 371516 334432 371568 334484
rect 440332 334432 440384 334484
rect 216588 334364 216640 334416
rect 300492 334364 300544 334416
rect 223488 334296 223540 334348
rect 303620 334296 303672 334348
rect 205548 333888 205600 333940
rect 296444 333888 296496 333940
rect 374644 333888 374696 333940
rect 445760 333888 445812 333940
rect 198648 333820 198700 333872
rect 295800 333820 295852 333872
rect 373816 333820 373868 333872
rect 448612 333820 448664 333872
rect 177948 333752 178000 333804
rect 288440 333752 288492 333804
rect 375012 333752 375064 333804
rect 452660 333752 452712 333804
rect 162768 333684 162820 333736
rect 284852 333684 284904 333736
rect 377404 333684 377456 333736
rect 459560 333684 459612 333736
rect 158628 333616 158680 333668
rect 282644 333616 282696 333668
rect 380532 333616 380584 333668
rect 470600 333616 470652 333668
rect 151728 333548 151780 333600
rect 281448 333548 281500 333600
rect 387616 333548 387668 333600
rect 492680 333548 492732 333600
rect 104164 333480 104216 333532
rect 266360 333480 266412 333532
rect 390928 333480 390980 333532
rect 502984 333480 503036 333532
rect 93124 333412 93176 333464
rect 262956 333412 263008 333464
rect 394608 333412 394660 333464
rect 515404 333412 515456 333464
rect 88984 333344 89036 333396
rect 261944 333344 261996 333396
rect 399300 333344 399352 333396
rect 530584 333344 530636 333396
rect 84108 333276 84160 333328
rect 400128 333276 400180 333328
rect 533344 333276 533396 333328
rect 39304 333208 39356 333260
rect 241796 333208 241848 333260
rect 401508 333208 401560 333260
rect 538220 333208 538272 333260
rect 209688 333140 209740 333192
rect 299112 333140 299164 333192
rect 227628 333072 227680 333124
rect 304632 333072 304684 333124
rect 260380 333004 260432 333056
rect 219256 332528 219308 332580
rect 302608 332528 302660 332580
rect 188988 332460 189040 332512
rect 291568 332460 291620 332512
rect 182088 332392 182140 332444
rect 290832 332392 290884 332444
rect 175188 332324 175240 332376
rect 288532 332324 288584 332376
rect 376208 332324 376260 332376
rect 456892 332324 456944 332376
rect 171048 332256 171100 332308
rect 287428 332256 287480 332308
rect 378508 332256 378560 332308
rect 463700 332256 463752 332308
rect 143448 332188 143500 332240
rect 274456 332188 274508 332240
rect 379428 332188 379480 332240
rect 466460 332188 466512 332240
rect 124128 332120 124180 332172
rect 271788 332120 271840 332172
rect 382832 332120 382884 332172
rect 477500 332120 477552 332172
rect 106188 332052 106240 332104
rect 267372 332052 267424 332104
rect 385316 332052 385368 332104
rect 485780 332052 485832 332104
rect 99288 331984 99340 332036
rect 264888 331984 264940 332036
rect 386328 331984 386380 332036
rect 489184 331984 489236 332036
rect 95148 331916 95200 331968
rect 264060 331916 264112 331968
rect 388720 331916 388772 331968
rect 496820 331916 496872 331968
rect 68284 331848 68336 331900
rect 250168 331848 250220 331900
rect 391848 331848 391900 331900
rect 506480 331848 506532 331900
rect 410616 331100 410668 331152
rect 411168 331100 411220 331152
rect 153108 330964 153160 331016
rect 282000 330964 282052 331016
rect 146208 330896 146260 330948
rect 277860 330896 277912 330948
rect 117228 330828 117280 330880
rect 270868 330828 270920 330880
rect 399668 330828 399720 330880
rect 485044 330828 485096 330880
rect 113088 330760 113140 330812
rect 269580 330760 269632 330812
rect 331588 330760 331640 330812
rect 389824 330760 389876 330812
rect 499580 330760 499632 330812
rect 111064 330692 111116 330744
rect 268476 330692 268528 330744
rect 81348 330624 81400 330676
rect 259644 330624 259696 330676
rect 392860 330692 392912 330744
rect 510620 330692 510672 330744
rect 394148 330624 394200 330676
rect 514760 330624 514812 330676
rect 61384 330556 61436 330608
rect 252560 330556 252612 330608
rect 331588 330556 331640 330608
rect 395160 330556 395212 330608
rect 517520 330556 517572 330608
rect 33784 330488 33836 330540
rect 234804 330420 234856 330472
rect 235264 330420 235316 330472
rect 236092 330420 236144 330472
rect 237012 330420 237064 330472
rect 237380 330420 237432 330472
rect 238484 330420 238536 330472
rect 241612 330488 241664 330540
rect 242532 330488 242584 330540
rect 244372 330488 244424 330540
rect 245108 330488 245160 330540
rect 247132 330488 247184 330540
rect 247316 330488 247368 330540
rect 248512 330488 248564 330540
rect 249432 330488 249484 330540
rect 249984 330488 250036 330540
rect 250904 330488 250956 330540
rect 251272 330488 251324 330540
rect 252008 330488 252060 330540
rect 253940 330488 253992 330540
rect 254584 330488 254636 330540
rect 255320 330488 255372 330540
rect 255688 330488 255740 330540
rect 258172 330488 258224 330540
rect 259000 330488 259052 330540
rect 265164 330488 265216 330540
rect 265900 330488 265952 330540
rect 266452 330488 266504 330540
rect 267004 330488 267056 330540
rect 270592 330488 270644 330540
rect 271328 330488 271380 330540
rect 271972 330488 272024 330540
rect 272432 330488 272484 330540
rect 285772 330488 285824 330540
rect 286324 330488 286376 330540
rect 287152 330488 287204 330540
rect 288164 330488 288216 330540
rect 291292 330488 291344 330540
rect 291844 330488 291896 330540
rect 294144 330488 294196 330540
rect 295156 330488 295208 330540
rect 299572 330488 299624 330540
rect 300584 330488 300636 330540
rect 300952 330488 301004 330540
rect 301688 330488 301740 330540
rect 311992 330488 312044 330540
rect 312636 330488 312688 330540
rect 313280 330488 313332 330540
rect 314108 330488 314160 330540
rect 317604 330488 317656 330540
rect 318524 330488 318576 330540
rect 318892 330488 318944 330540
rect 319536 330488 319588 330540
rect 320180 330488 320232 330540
rect 321008 330488 321060 330540
rect 321652 330488 321704 330540
rect 322112 330488 322164 330540
rect 323124 330488 323176 330540
rect 323952 330488 324004 330540
rect 324320 330488 324372 330540
rect 324688 330488 324740 330540
rect 325792 330488 325844 330540
rect 326528 330488 326580 330540
rect 329932 330488 329984 330540
rect 330944 330488 330996 330540
rect 331496 330488 331548 330540
rect 331956 330488 332008 330540
rect 332600 330488 332652 330540
rect 333428 330488 333480 330540
rect 334072 330488 334124 330540
rect 334532 330488 334584 330540
rect 335452 330488 335504 330540
rect 336372 330488 336424 330540
rect 338120 330488 338172 330540
rect 338580 330488 338632 330540
rect 349988 330488 350040 330540
rect 350448 330488 350500 330540
rect 362408 330488 362460 330540
rect 362868 330488 362920 330540
rect 381360 330488 381412 330540
rect 382096 330488 382148 330540
rect 396356 330488 396408 330540
rect 519544 330488 519596 330540
rect 244464 330420 244516 330472
rect 254032 330420 254084 330472
rect 254952 330420 255004 330472
rect 255412 330420 255464 330472
rect 256056 330420 256108 330472
rect 324412 330420 324464 330472
rect 325424 330420 325476 330472
rect 331312 330420 331364 330472
rect 332324 330420 332376 330472
rect 338212 330420 338264 330472
rect 338948 330420 339000 330472
rect 414296 330420 414348 330472
rect 415124 330420 415176 330472
rect 119988 329332 120040 329384
rect 269120 329332 269172 329384
rect 58624 329264 58676 329316
rect 248696 329264 248748 329316
rect 47584 329196 47636 329248
rect 246580 329196 246632 329248
rect 32404 329128 32456 329180
rect 240324 329128 240376 329180
rect 397368 329128 397420 329180
rect 524420 329128 524472 329180
rect 36544 329060 36596 329112
rect 245660 329060 245712 329112
rect 400772 329060 400824 329112
rect 535460 329060 535512 329112
rect 329840 328040 329892 328092
rect 330576 328040 330628 328092
rect 14464 327700 14516 327752
rect 237748 327700 237800 327752
rect 314752 327156 314804 327208
rect 315580 327156 315632 327208
rect 276204 326408 276256 326460
rect 302516 326451 302568 326460
rect 302516 326417 302525 326451
rect 302525 326417 302559 326451
rect 302559 326417 302568 326451
rect 302516 326408 302568 326417
rect 309232 326408 309284 326460
rect 310060 326408 310112 326460
rect 274732 326340 274784 326392
rect 275744 326340 275796 326392
rect 234712 326272 234764 326324
rect 235540 326272 235592 326324
rect 277492 326340 277544 326392
rect 277676 326340 277728 326392
rect 280252 326340 280304 326392
rect 280896 326340 280948 326392
rect 302332 326340 302384 326392
rect 303160 326340 303212 326392
rect 305000 326340 305052 326392
rect 305368 326340 305420 326392
rect 306380 326340 306432 326392
rect 307484 326340 307536 326392
rect 307760 326340 307812 326392
rect 308588 326340 308640 326392
rect 309140 326340 309192 326392
rect 309692 326340 309744 326392
rect 310612 326340 310664 326392
rect 311164 326340 311216 326392
rect 276204 326204 276256 326256
rect 277492 326204 277544 326256
rect 278320 326204 278372 326256
rect 305092 326204 305144 326256
rect 305736 326204 305788 326256
rect 305184 326136 305236 326188
rect 306104 326136 306156 326188
rect 421656 325592 421708 325644
rect 579896 325592 579948 325644
rect 302516 323595 302568 323604
rect 302516 323561 302525 323595
rect 302525 323561 302559 323595
rect 302559 323561 302568 323595
rect 302516 323552 302568 323561
rect 276112 321512 276164 321564
rect 276296 321512 276348 321564
rect 555424 313216 555476 313268
rect 580172 313216 580224 313268
rect 3332 215228 3384 215280
rect 232596 215228 232648 215280
rect 3424 45500 3476 45552
rect 226984 45500 227036 45552
rect 3424 20612 3476 20664
rect 414940 20612 414992 20664
rect 431224 20612 431276 20664
rect 579988 20612 580040 20664
rect 157248 18572 157300 18624
rect 282184 18572 282236 18624
rect 161296 17212 161348 17264
rect 284392 17212 284444 17264
rect 139308 15852 139360 15904
rect 277584 15852 277636 15904
rect 252376 14424 252428 14476
rect 311992 14424 312044 14476
rect 184940 13336 184992 13388
rect 291292 13336 291344 13388
rect 125876 13268 125928 13320
rect 233976 13268 234028 13320
rect 164148 13200 164200 13252
rect 284484 13200 284536 13252
rect 149980 13132 150032 13184
rect 280252 13132 280304 13184
rect 128176 13064 128228 13116
rect 273444 13064 273496 13116
rect 212172 12180 212224 12232
rect 233884 12180 233936 12232
rect 182548 12112 182600 12164
rect 224224 12112 224276 12164
rect 175924 12044 175976 12096
rect 228364 12044 228416 12096
rect 164884 11976 164936 12028
rect 231124 11976 231176 12028
rect 154212 11908 154264 11960
rect 232504 11908 232556 11960
rect 251088 11908 251140 11960
rect 291844 11908 291896 11960
rect 167644 11840 167696 11892
rect 285772 11840 285824 11892
rect 78588 11772 78640 11824
rect 258356 11772 258408 11824
rect 74448 11704 74500 11756
rect 256884 11704 256936 11756
rect 440332 11704 440384 11756
rect 441528 11704 441580 11756
rect 448612 11704 448664 11756
rect 449808 11704 449860 11756
rect 160100 11636 160152 11688
rect 161296 11636 161348 11688
rect 95056 10956 95108 11008
rect 263692 10956 263744 11008
rect 428464 10956 428516 11008
rect 430856 10956 430908 11008
rect 91008 10888 91060 10940
rect 262404 10888 262456 10940
rect 70308 10820 70360 10872
rect 255596 10820 255648 10872
rect 67548 10752 67600 10804
rect 255504 10752 255556 10804
rect 63224 10684 63276 10736
rect 254216 10684 254268 10736
rect 60648 10616 60700 10668
rect 252744 10616 252796 10668
rect 260656 10616 260708 10668
rect 286324 10616 286376 10668
rect 56508 10548 56560 10600
rect 251272 10548 251324 10600
rect 253848 10548 253900 10600
rect 289084 10548 289136 10600
rect 53748 10480 53800 10532
rect 249984 10480 250036 10532
rect 271788 10480 271840 10532
rect 317604 10480 317656 10532
rect 49608 10412 49660 10464
rect 249892 10412 249944 10464
rect 269028 10412 269080 10464
rect 317512 10412 317564 10464
rect 45468 10344 45520 10396
rect 248604 10344 248656 10396
rect 264888 10344 264940 10396
rect 316132 10344 316184 10396
rect 41328 10276 41380 10328
rect 247132 10276 247184 10328
rect 256608 10276 256660 10328
rect 313464 10276 313516 10328
rect 357164 10276 357216 10328
rect 392584 10276 392636 10328
rect 97908 10208 97960 10260
rect 265072 10208 265124 10260
rect 102048 10140 102100 10192
rect 265164 10140 265216 10192
rect 104532 10072 104584 10124
rect 266452 10072 266504 10124
rect 108948 10004 109000 10056
rect 267832 10004 267884 10056
rect 111616 9936 111668 9988
rect 269304 9936 269356 9988
rect 115848 9868 115900 9920
rect 270684 9868 270736 9920
rect 119804 9800 119856 9852
rect 270592 9800 270644 9852
rect 122748 9732 122800 9784
rect 271972 9732 272024 9784
rect 209780 9596 209832 9648
rect 299664 9596 299716 9648
rect 417516 9596 417568 9648
rect 420184 9596 420236 9648
rect 206192 9528 206244 9580
rect 298192 9528 298244 9580
rect 202696 9460 202748 9512
rect 296812 9460 296864 9512
rect 199108 9392 199160 9444
rect 295524 9392 295576 9444
rect 195612 9324 195664 9376
rect 294144 9324 294196 9376
rect 192024 9256 192076 9308
rect 294052 9256 294104 9308
rect 135260 9188 135312 9240
rect 276112 9188 276164 9240
rect 131764 9120 131816 9172
rect 274916 9120 274968 9172
rect 37188 9052 37240 9104
rect 245936 9052 245988 9104
rect 248788 9052 248840 9104
rect 310796 9052 310848 9104
rect 418804 9052 418856 9104
rect 427268 9052 427320 9104
rect 33600 8984 33652 9036
rect 244372 8984 244424 9036
rect 245200 8984 245252 9036
rect 310704 8984 310756 9036
rect 353944 8984 353996 9036
rect 370596 8984 370648 9036
rect 372436 8984 372488 9036
rect 445024 8984 445076 9036
rect 8760 8916 8812 8968
rect 237472 8916 237524 8968
rect 238116 8916 238168 8968
rect 307944 8916 307996 8968
rect 353024 8916 353076 8968
rect 382372 8916 382424 8968
rect 382924 8916 382976 8968
rect 416688 8916 416740 8968
rect 417424 8916 417476 8968
rect 494704 8916 494756 8968
rect 126980 8848 127032 8900
rect 213184 8848 213236 8900
rect 213368 8848 213420 8900
rect 299572 8848 299624 8900
rect 216864 8780 216916 8832
rect 300952 8780 301004 8832
rect 220452 8712 220504 8764
rect 302424 8712 302476 8764
rect 223948 8644 224000 8696
rect 303712 8644 303764 8696
rect 227536 8576 227588 8628
rect 305276 8576 305328 8628
rect 231032 8508 231084 8560
rect 305184 8508 305236 8560
rect 234988 8440 235040 8492
rect 306656 8440 306708 8492
rect 241704 8372 241756 8424
rect 309416 8372 309468 8424
rect 421564 8304 421616 8356
rect 423772 8304 423824 8356
rect 137652 8236 137704 8288
rect 277676 8236 277728 8288
rect 372344 8236 372396 8288
rect 442632 8236 442684 8288
rect 134156 8168 134208 8220
rect 276204 8168 276256 8220
rect 403992 8168 404044 8220
rect 545488 8168 545540 8220
rect 79692 8100 79744 8152
rect 76196 8032 76248 8084
rect 258356 8100 258408 8152
rect 259552 8100 259604 8152
rect 265348 8100 265400 8152
rect 316224 8100 316276 8152
rect 405372 8100 405424 8152
rect 549076 8100 549128 8152
rect 258264 8032 258316 8084
rect 72608 7964 72660 8016
rect 256792 7964 256844 8016
rect 261760 8032 261812 8084
rect 314752 8032 314804 8084
rect 405464 8032 405516 8084
rect 552664 8032 552716 8084
rect 30104 7896 30156 7948
rect 243084 7896 243136 7948
rect 251180 7896 251232 7948
rect 314844 7964 314896 8016
rect 406752 7964 406804 8016
rect 556160 7964 556212 8016
rect 26516 7828 26568 7880
rect 242992 7828 243044 7880
rect 254676 7828 254728 7880
rect 313372 7896 313424 7948
rect 408224 7896 408276 7948
rect 559748 7896 559800 7948
rect 312084 7828 312136 7880
rect 409512 7828 409564 7880
rect 563244 7828 563296 7880
rect 21824 7760 21876 7812
rect 241796 7760 241848 7812
rect 247592 7760 247644 7812
rect 310612 7760 310664 7812
rect 410984 7760 411036 7812
rect 566832 7760 566884 7812
rect 17040 7692 17092 7744
rect 240140 7692 240192 7744
rect 244096 7692 244148 7744
rect 309232 7692 309284 7744
rect 410892 7692 410944 7744
rect 570328 7692 570380 7744
rect 12348 7624 12400 7676
rect 237380 7624 237432 7676
rect 240508 7624 240560 7676
rect 309324 7624 309376 7676
rect 412272 7624 412324 7676
rect 573916 7624 573968 7676
rect 4068 7556 4120 7608
rect 236184 7556 236236 7608
rect 237012 7556 237064 7608
rect 307852 7556 307904 7608
rect 413744 7556 413796 7608
rect 577412 7556 577464 7608
rect 141240 7488 141292 7540
rect 277492 7488 277544 7540
rect 371056 7488 371108 7540
rect 144736 7420 144788 7472
rect 278964 7420 279016 7472
rect 369676 7420 369728 7472
rect 148324 7352 148376 7404
rect 280344 7352 280396 7404
rect 368388 7352 368440 7404
rect 432052 7352 432104 7404
rect 151820 7284 151872 7336
rect 281724 7284 281776 7336
rect 368296 7284 368348 7336
rect 428464 7284 428516 7336
rect 432604 7488 432656 7540
rect 434444 7488 434496 7540
rect 435364 7488 435416 7540
rect 437940 7488 437992 7540
rect 439136 7352 439188 7404
rect 435548 7284 435600 7336
rect 155408 7216 155460 7268
rect 283012 7216 283064 7268
rect 367008 7216 367060 7268
rect 424968 7216 425020 7268
rect 158904 7148 158956 7200
rect 283104 7148 283156 7200
rect 365536 7148 365588 7200
rect 421380 7148 421432 7200
rect 229836 7080 229888 7132
rect 305092 7080 305144 7132
rect 364156 7080 364208 7132
rect 417884 7080 417936 7132
rect 233424 7012 233476 7064
rect 306564 7012 306616 7064
rect 362592 7012 362644 7064
rect 414296 7012 414348 7064
rect 234620 6808 234672 6860
rect 580172 6808 580224 6860
rect 169576 6740 169628 6792
rect 287244 6740 287296 6792
rect 382004 6740 382056 6792
rect 476948 6740 477000 6792
rect 166080 6672 166132 6724
rect 285864 6672 285916 6724
rect 384856 6672 384908 6724
rect 481732 6672 481784 6724
rect 130568 6604 130620 6656
rect 274824 6604 274876 6656
rect 384764 6604 384816 6656
rect 485228 6604 485280 6656
rect 69112 6536 69164 6588
rect 255412 6536 255464 6588
rect 386328 6536 386380 6588
rect 488816 6536 488868 6588
rect 65524 6468 65576 6520
rect 254032 6468 254084 6520
rect 387708 6468 387760 6520
rect 492312 6468 492364 6520
rect 62028 6400 62080 6452
rect 254124 6400 254176 6452
rect 389088 6400 389140 6452
rect 495900 6400 495952 6452
rect 58440 6332 58492 6384
rect 252652 6332 252704 6384
rect 299664 6332 299716 6384
rect 316684 6332 316736 6384
rect 390192 6332 390244 6384
rect 499396 6332 499448 6384
rect 54944 6264 54996 6316
rect 251364 6264 251416 6316
rect 259460 6264 259512 6316
rect 295984 6264 296036 6316
rect 303160 6264 303212 6316
rect 327724 6264 327776 6316
rect 390376 6264 390428 6316
rect 502892 6264 502944 6316
rect 51356 6196 51408 6248
rect 250076 6196 250128 6248
rect 268844 6196 268896 6248
rect 317696 6196 317748 6248
rect 371884 6196 371936 6248
rect 378876 6196 378928 6248
rect 391664 6196 391716 6248
rect 506480 6196 506532 6248
rect 47860 6128 47912 6180
rect 248512 6128 248564 6180
rect 257068 6128 257120 6180
rect 313280 6128 313332 6180
rect 370504 6128 370556 6180
rect 385960 6128 386012 6180
rect 393136 6128 393188 6180
rect 510068 6128 510120 6180
rect 173164 6060 173216 6112
rect 287152 6060 287204 6112
rect 382096 6060 382148 6112
rect 473452 6060 473504 6112
rect 176660 5992 176712 6044
rect 288624 5992 288676 6044
rect 380716 5992 380768 6044
rect 469864 5992 469916 6044
rect 180248 5924 180300 5976
rect 290004 5924 290056 5976
rect 379428 5924 379480 5976
rect 466276 5924 466328 5976
rect 468484 5924 468536 5976
rect 474556 5924 474608 5976
rect 183744 5856 183796 5908
rect 291384 5856 291436 5908
rect 377956 5856 378008 5908
rect 462780 5856 462832 5908
rect 187332 5788 187384 5840
rect 292672 5788 292724 5840
rect 377864 5788 377916 5840
rect 459192 5788 459244 5840
rect 190828 5720 190880 5772
rect 292764 5720 292816 5772
rect 376668 5720 376720 5772
rect 455696 5720 455748 5772
rect 194416 5652 194468 5704
rect 294236 5652 294288 5704
rect 375196 5652 375248 5704
rect 452108 5652 452160 5704
rect 363604 5516 363656 5568
rect 367008 5516 367060 5568
rect 475384 5516 475436 5568
rect 480536 5516 480588 5568
rect 486424 5516 486476 5568
rect 487620 5516 487672 5568
rect 497464 5516 497516 5568
rect 498200 5516 498252 5568
rect 504364 5516 504416 5568
rect 505376 5516 505428 5568
rect 186136 5448 186188 5500
rect 215944 5448 215996 5500
rect 218060 5448 218112 5500
rect 302516 5448 302568 5500
rect 355876 5448 355928 5500
rect 391848 5448 391900 5500
rect 402704 5448 402756 5500
rect 540796 5448 540848 5500
rect 189724 5380 189776 5432
rect 214288 5380 214340 5432
rect 214472 5380 214524 5432
rect 301044 5380 301096 5432
rect 357256 5380 357308 5432
rect 395252 5380 395304 5432
rect 404176 5380 404228 5432
rect 544384 5380 544436 5432
rect 210976 5312 211028 5364
rect 299756 5312 299808 5364
rect 358636 5312 358688 5364
rect 400128 5312 400180 5364
rect 404084 5312 404136 5364
rect 547880 5312 547932 5364
rect 136456 5244 136508 5296
rect 204904 5244 204956 5296
rect 207388 5244 207440 5296
rect 298284 5244 298336 5296
rect 358544 5244 358596 5296
rect 398932 5244 398984 5296
rect 405556 5244 405608 5296
rect 551468 5244 551520 5296
rect 203892 5176 203944 5228
rect 296904 5176 296956 5228
rect 359924 5176 359976 5228
rect 402520 5176 402572 5228
rect 406844 5176 406896 5228
rect 554964 5176 555016 5228
rect 132960 5108 133012 5160
rect 274732 5108 274784 5160
rect 278320 5108 278372 5160
rect 320364 5108 320416 5160
rect 359832 5108 359884 5160
rect 403624 5108 403676 5160
rect 408316 5108 408368 5160
rect 558552 5108 558604 5160
rect 129372 5040 129424 5092
rect 274640 5040 274692 5092
rect 274824 5040 274876 5092
rect 318892 5040 318944 5092
rect 361304 5040 361356 5092
rect 406016 5040 406068 5092
rect 409604 5040 409656 5092
rect 562048 5040 562100 5092
rect 7656 4972 7708 5024
rect 236092 4972 236144 5024
rect 246396 4972 246448 5024
rect 310520 4972 310572 5024
rect 361396 4972 361448 5024
rect 407212 4972 407264 5024
rect 409696 4972 409748 5024
rect 565636 4972 565688 5024
rect 2872 4904 2924 4956
rect 234712 4904 234764 4956
rect 242900 4904 242952 4956
rect 309140 4904 309192 4956
rect 362684 4904 362736 4956
rect 410800 4904 410852 4956
rect 411076 4904 411128 4956
rect 569132 4904 569184 4956
rect 1676 4836 1728 4888
rect 234804 4836 234856 4888
rect 239312 4836 239364 4888
rect 307760 4836 307812 4888
rect 361212 4836 361264 4888
rect 409604 4836 409656 4888
rect 412364 4836 412416 4888
rect 572720 4836 572772 4888
rect 572 4768 624 4820
rect 234896 4768 234948 4820
rect 235816 4768 235868 4820
rect 306380 4768 306432 4820
rect 362776 4768 362828 4820
rect 413100 4768 413152 4820
rect 413836 4768 413888 4820
rect 576308 4768 576360 4820
rect 193220 4700 193272 4752
rect 220084 4700 220136 4752
rect 221556 4700 221608 4752
rect 302332 4700 302384 4752
rect 355784 4700 355836 4752
rect 388260 4700 388312 4752
rect 401324 4700 401376 4752
rect 537208 4700 537260 4752
rect 171968 4632 172020 4684
rect 222844 4632 222896 4684
rect 225144 4632 225196 4684
rect 303804 4632 303856 4684
rect 354496 4632 354548 4684
rect 384764 4632 384816 4684
rect 399852 4632 399904 4684
rect 533712 4632 533764 4684
rect 228732 4564 228784 4616
rect 305000 4564 305052 4616
rect 353116 4564 353168 4616
rect 381176 4564 381228 4616
rect 398656 4564 398708 4616
rect 530124 4564 530176 4616
rect 232228 4496 232280 4548
rect 306472 4496 306524 4548
rect 351736 4496 351788 4548
rect 377680 4496 377732 4548
rect 398564 4496 398616 4548
rect 526628 4496 526680 4548
rect 281908 4428 281960 4480
rect 321744 4428 321796 4480
rect 350264 4428 350316 4480
rect 374092 4428 374144 4480
rect 397092 4428 397144 4480
rect 523040 4428 523092 4480
rect 285404 4360 285456 4412
rect 323032 4360 323084 4412
rect 395804 4360 395856 4412
rect 519544 4360 519596 4412
rect 288992 4292 289044 4344
rect 323124 4292 323176 4344
rect 394424 4292 394476 4344
rect 515956 4292 516008 4344
rect 200304 4224 200356 4276
rect 208952 4224 209004 4276
rect 292580 4224 292632 4276
rect 324596 4224 324648 4276
rect 392952 4224 393004 4276
rect 512460 4224 512512 4276
rect 11152 4088 11204 4140
rect 18604 4088 18656 4140
rect 34796 4088 34848 4140
rect 36544 4088 36596 4140
rect 78496 4088 78548 4140
rect 82084 4020 82136 4072
rect 143540 4156 143592 4208
rect 144828 4156 144880 4208
rect 168380 4156 168432 4208
rect 169668 4156 169720 4208
rect 201500 4156 201552 4208
rect 202788 4156 202840 4208
rect 226340 4156 226392 4208
rect 227628 4156 227680 4208
rect 388444 4156 388496 4208
rect 389456 4156 389508 4208
rect 395344 4156 395396 4208
rect 396540 4156 396592 4208
rect 259736 4088 259788 4140
rect 309048 4088 309100 4140
rect 330116 4088 330168 4140
rect 332692 4088 332744 4140
rect 336004 4088 336056 4140
rect 343456 4088 343508 4140
rect 350448 4088 350500 4140
rect 351828 4088 351880 4140
rect 375288 4088 375340 4140
rect 402612 4088 402664 4140
rect 258172 4020 258224 4072
rect 307944 4020 307996 4072
rect 330024 4020 330076 4072
rect 343548 4020 343600 4072
rect 348056 4020 348108 4072
rect 350356 4020 350408 4072
rect 372896 4020 372948 4072
rect 402796 4020 402848 4072
rect 543188 4020 543240 4072
rect 43076 3952 43128 4004
rect 51724 3952 51776 4004
rect 53656 3952 53708 4004
rect 57244 3952 57296 4004
rect 75000 3952 75052 4004
rect 258080 3952 258132 4004
rect 305552 3952 305604 4004
rect 328552 3952 328604 4004
rect 329196 3952 329248 4004
rect 335452 3952 335504 4004
rect 343364 3952 343416 4004
rect 349252 3952 349304 4004
rect 353208 3952 353260 4004
rect 379980 3952 380032 4004
rect 404268 3952 404320 4004
rect 546684 3952 546736 4004
rect 38384 3884 38436 3936
rect 47584 3884 47636 3936
rect 50160 3884 50212 3936
rect 68284 3884 68336 3936
rect 71504 3884 71556 3936
rect 256700 3884 256752 3936
rect 301964 3884 302016 3936
rect 5264 3816 5316 3868
rect 7564 3816 7616 3868
rect 41880 3816 41932 3868
rect 54484 3816 54536 3868
rect 67916 3816 67968 3868
rect 255320 3816 255372 3868
rect 297272 3816 297324 3868
rect 325792 3884 325844 3936
rect 320916 3816 320968 3868
rect 35992 3748 36044 3800
rect 50344 3748 50396 3800
rect 64328 3748 64380 3800
rect 253940 3748 253992 3800
rect 293684 3748 293736 3800
rect 324320 3748 324372 3800
rect 324412 3748 324464 3800
rect 334256 3884 334308 3936
rect 344284 3884 344336 3936
rect 351644 3884 351696 3936
rect 354588 3884 354640 3936
rect 387156 3884 387208 3936
rect 405648 3884 405700 3936
rect 550272 3884 550324 3936
rect 329104 3816 329156 3868
rect 333888 3816 333940 3868
rect 336924 3816 336976 3868
rect 345756 3816 345808 3868
rect 356336 3816 356388 3868
rect 357348 3816 357400 3868
rect 23020 3680 23072 3732
rect 39304 3680 39356 3732
rect 20628 3612 20680 3664
rect 43444 3680 43496 3732
rect 45376 3680 45428 3732
rect 58624 3680 58676 3732
rect 60832 3680 60884 3732
rect 252836 3680 252888 3732
rect 291384 3680 291436 3732
rect 327264 3748 327316 3800
rect 331220 3748 331272 3800
rect 331496 3748 331548 3800
rect 346308 3748 346360 3800
rect 326804 3680 326856 3732
rect 335636 3680 335688 3732
rect 347596 3680 347648 3732
rect 39580 3612 39632 3664
rect 18236 3544 18288 3596
rect 28908 3544 28960 3596
rect 35164 3544 35216 3596
rect 40684 3544 40736 3596
rect 41328 3544 41380 3596
rect 48964 3544 49016 3596
rect 49608 3544 49660 3596
rect 52552 3544 52604 3596
rect 53748 3544 53800 3596
rect 248696 3612 248748 3664
rect 286600 3612 286652 3664
rect 323216 3612 323268 3664
rect 247224 3544 247276 3596
rect 279516 3544 279568 3596
rect 32312 3476 32364 3528
rect 32404 3476 32456 3528
rect 244464 3476 244516 3528
rect 249984 3476 250036 3528
rect 251088 3476 251140 3528
rect 255872 3476 255924 3528
rect 256608 3476 256660 3528
rect 262956 3476 263008 3528
rect 263508 3476 263560 3528
rect 264152 3476 264204 3528
rect 264888 3476 264940 3528
rect 266544 3476 266596 3528
rect 267648 3476 267700 3528
rect 267740 3476 267792 3528
rect 269028 3476 269080 3528
rect 271236 3476 271288 3528
rect 271788 3476 271840 3528
rect 273628 3476 273680 3528
rect 274548 3476 274600 3528
rect 280712 3476 280764 3528
rect 281448 3476 281500 3528
rect 284300 3544 284352 3596
rect 321836 3544 321888 3596
rect 324228 3612 324280 3664
rect 325608 3612 325660 3664
rect 335544 3612 335596 3664
rect 347136 3612 347188 3664
rect 358728 3748 358780 3800
rect 390652 3816 390704 3868
rect 407028 3816 407080 3868
rect 553768 3816 553820 3868
rect 358084 3680 358136 3732
rect 363512 3680 363564 3732
rect 394240 3748 394292 3800
rect 406936 3748 406988 3800
rect 557356 3748 557408 3800
rect 397736 3680 397788 3732
rect 408408 3680 408460 3732
rect 560852 3680 560904 3732
rect 320180 3476 320232 3528
rect 323400 3544 323452 3596
rect 334072 3544 334124 3596
rect 342076 3544 342128 3596
rect 346952 3544 347004 3596
rect 347688 3544 347740 3596
rect 358728 3612 358780 3664
rect 360016 3612 360068 3664
rect 401324 3612 401376 3664
rect 409788 3612 409840 3664
rect 564440 3612 564492 3664
rect 322112 3476 322164 3528
rect 331588 3476 331640 3528
rect 332508 3476 332560 3528
rect 336280 3476 336332 3528
rect 338120 3476 338172 3528
rect 345664 3476 345716 3528
rect 352840 3476 352892 3528
rect 359924 3544 359976 3596
rect 360108 3544 360160 3596
rect 404820 3544 404872 3596
rect 411168 3544 411220 3596
rect 568028 3544 568080 3596
rect 361120 3476 361172 3528
rect 361488 3476 361540 3528
rect 408408 3476 408460 3528
rect 412456 3476 412508 3528
rect 571524 3476 571576 3528
rect 13544 3408 13596 3460
rect 22744 3408 22796 3460
rect 25320 3408 25372 3460
rect 241612 3408 241664 3460
rect 272432 3408 272484 3460
rect 318984 3408 319036 3460
rect 319720 3408 319772 3460
rect 332600 3408 332652 3460
rect 335084 3408 335136 3460
rect 338304 3408 338356 3460
rect 348976 3408 349028 3460
rect 362316 3408 362368 3460
rect 362868 3408 362920 3460
rect 411904 3408 411956 3460
rect 412548 3408 412600 3460
rect 575112 3408 575164 3460
rect 19432 3340 19484 3392
rect 25504 3340 25556 3392
rect 31300 3340 31352 3392
rect 33784 3340 33836 3392
rect 44272 3340 44324 3392
rect 45468 3340 45520 3392
rect 46664 3340 46716 3392
rect 56048 3340 56100 3392
rect 56508 3340 56560 3392
rect 59636 3340 59688 3392
rect 60648 3340 60700 3392
rect 66720 3340 66772 3392
rect 67548 3340 67600 3392
rect 77392 3340 77444 3392
rect 78588 3340 78640 3392
rect 80888 3340 80940 3392
rect 81348 3340 81400 3392
rect 83280 3340 83332 3392
rect 84108 3340 84160 3392
rect 84476 3340 84528 3392
rect 87604 3340 87656 3392
rect 87972 3340 88024 3392
rect 88984 3340 89036 3392
rect 90364 3340 90416 3392
rect 91008 3340 91060 3392
rect 91560 3340 91612 3392
rect 93124 3340 93176 3392
rect 85672 3272 85724 3324
rect 261024 3340 261076 3392
rect 287796 3340 287848 3392
rect 288348 3340 288400 3392
rect 298468 3340 298520 3392
rect 299388 3340 299440 3392
rect 304356 3340 304408 3392
rect 304908 3340 304960 3392
rect 306748 3340 306800 3392
rect 328736 3340 328788 3392
rect 334164 3340 334216 3392
rect 348516 3340 348568 3392
rect 355232 3340 355284 3392
rect 97448 3272 97500 3324
rect 97908 3272 97960 3324
rect 98644 3272 98696 3324
rect 99288 3272 99340 3324
rect 101036 3272 101088 3324
rect 102048 3272 102100 3324
rect 262312 3272 262364 3324
rect 310244 3272 310296 3324
rect 329840 3272 329892 3324
rect 350540 3272 350592 3324
rect 371700 3340 371752 3392
rect 382188 3340 382240 3392
rect 475752 3340 475804 3392
rect 489184 3340 489236 3392
rect 489920 3340 489972 3392
rect 369400 3272 369452 3324
rect 380624 3272 380676 3324
rect 468668 3272 468720 3324
rect 485044 3272 485096 3324
rect 502984 3272 503036 3324
rect 504180 3272 504232 3324
rect 515404 3272 515456 3324
rect 517152 3272 517204 3324
rect 519636 3272 519688 3324
rect 521844 3272 521896 3324
rect 522304 3272 522356 3324
rect 524236 3272 524288 3324
rect 530584 3340 530636 3392
rect 531320 3340 531372 3392
rect 533344 3340 533396 3392
rect 534908 3340 534960 3392
rect 539600 3340 539652 3392
rect 540244 3340 540296 3392
rect 541992 3340 542044 3392
rect 532516 3272 532568 3324
rect 92756 3204 92808 3256
rect 262496 3204 262548 3256
rect 311440 3204 311492 3256
rect 329932 3204 329984 3256
rect 57244 3136 57296 3188
rect 61384 3136 61436 3188
rect 93952 3136 94004 3188
rect 95056 3136 95108 3188
rect 96252 3136 96304 3188
rect 263784 3136 263836 3188
rect 312636 3136 312688 3188
rect 331496 3204 331548 3256
rect 349068 3204 349120 3256
rect 365812 3204 365864 3256
rect 377772 3204 377824 3256
rect 461584 3204 461636 3256
rect 526444 3204 526496 3256
rect 527824 3204 527876 3256
rect 330392 3136 330444 3188
rect 333244 3136 333296 3188
rect 342168 3136 342220 3188
rect 344560 3136 344612 3188
rect 347044 3136 347096 3188
rect 354036 3136 354088 3188
rect 89168 3068 89220 3120
rect 102232 3068 102284 3120
rect 104164 3068 104216 3120
rect 105728 3068 105780 3120
rect 106188 3068 106240 3120
rect 106924 3068 106976 3120
rect 107568 3068 107620 3120
rect 108120 3068 108172 3120
rect 108948 3068 109000 3120
rect 109316 3068 109368 3120
rect 111064 3068 111116 3120
rect 265256 3068 265308 3120
rect 313832 3068 313884 3120
rect 331404 3068 331456 3120
rect 338672 3068 338724 3120
rect 339592 3068 339644 3120
rect 349804 3068 349856 3120
rect 357532 3068 357584 3120
rect 27712 3000 27764 3052
rect 29644 3000 29696 3052
rect 73804 3000 73856 3052
rect 74448 3000 74500 3052
rect 103336 3000 103388 3052
rect 266636 3000 266688 3052
rect 296076 3000 296128 3052
rect 296628 3000 296680 3052
rect 315028 3000 315080 3052
rect 331220 3000 331272 3052
rect 337476 3000 337528 3052
rect 338212 3000 338264 3052
rect 348424 3000 348476 3052
rect 364616 3136 364668 3188
rect 375104 3136 375156 3188
rect 454500 3136 454552 3188
rect 456800 3136 456852 3188
rect 458088 3136 458140 3188
rect 512644 3136 512696 3188
rect 513564 3136 513616 3188
rect 373908 3068 373960 3120
rect 447416 3068 447468 3120
rect 371148 3000 371200 3052
rect 440332 3000 440384 3052
rect 99840 2932 99892 2984
rect 9956 2864 10008 2916
rect 14464 2864 14516 2916
rect 110512 2932 110564 2984
rect 267924 2932 267976 2984
rect 317328 2932 317380 2984
rect 332784 2932 332836 2984
rect 355968 2932 356020 2984
rect 369768 2932 369820 2984
rect 433248 2932 433300 2984
rect 114008 2864 114060 2916
rect 114468 2864 114520 2916
rect 115204 2864 115256 2916
rect 115848 2864 115900 2916
rect 116400 2864 116452 2916
rect 117228 2864 117280 2916
rect 118792 2864 118844 2916
rect 119804 2864 119856 2916
rect 117596 2796 117648 2848
rect 270776 2864 270828 2916
rect 276020 2864 276072 2916
rect 277308 2864 277360 2916
rect 318524 2864 318576 2916
rect 332876 2864 332928 2916
rect 365628 2864 365680 2916
rect 422576 2864 422628 2916
rect 121092 2796 121144 2848
rect 272064 2796 272116 2848
rect 316224 2796 316276 2848
rect 331312 2796 331364 2848
rect 364248 2796 364300 2848
rect 415492 2796 415544 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 89364 703582 89668 703610
rect 8128 700330 8156 703520
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 24320 699718 24348 703520
rect 40512 700466 40540 703520
rect 40500 700460 40552 700466
rect 40500 700402 40552 700408
rect 41328 700460 41380 700466
rect 41328 700402 41380 700408
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3146 658200 3202 658209
rect 3146 658135 3202 658144
rect 3160 656946 3188 658135
rect 3148 656940 3200 656946
rect 3148 656882 3200 656888
rect 2962 619168 3018 619177
rect 2962 619103 3018 619112
rect 2976 618322 3004 619103
rect 2964 618316 3016 618322
rect 2964 618258 3016 618264
rect 3330 606112 3386 606121
rect 3330 606047 3386 606056
rect 3344 605878 3372 606047
rect 3332 605872 3384 605878
rect 3332 605814 3384 605820
rect 3330 566944 3386 566953
rect 3330 566879 3386 566888
rect 3344 565894 3372 566879
rect 3332 565888 3384 565894
rect 3332 565830 3384 565836
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 3330 514856 3386 514865
rect 3330 514791 3332 514800
rect 3384 514791 3386 514800
rect 3332 514762 3384 514768
rect 3238 501800 3294 501809
rect 3238 501735 3294 501744
rect 3252 501022 3280 501735
rect 3240 501016 3292 501022
rect 3240 500958 3292 500964
rect 3436 460562 3464 684247
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 465746 3556 671191
rect 3606 632088 3662 632097
rect 3606 632023 3662 632032
rect 3620 465882 3648 632023
rect 3698 580000 3754 580009
rect 3698 579935 3754 579944
rect 3712 466018 3740 579935
rect 3790 527912 3846 527921
rect 3790 527847 3846 527856
rect 3804 466154 3832 527847
rect 3974 475688 4030 475697
rect 3974 475623 4030 475632
rect 3804 466126 3924 466154
rect 3712 465990 3832 466018
rect 3620 465854 3740 465882
rect 3528 465718 3648 465746
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3528 462398 3556 462567
rect 3516 462392 3568 462398
rect 3516 462334 3568 462340
rect 3424 460556 3476 460562
rect 3424 460498 3476 460504
rect 3620 460494 3648 465718
rect 3608 460488 3660 460494
rect 3608 460430 3660 460436
rect 3712 460426 3740 465854
rect 3700 460420 3752 460426
rect 3700 460362 3752 460368
rect 3804 460358 3832 465990
rect 3792 460352 3844 460358
rect 3792 460294 3844 460300
rect 3896 460290 3924 466126
rect 3884 460284 3936 460290
rect 3884 460226 3936 460232
rect 3988 460222 4016 475623
rect 24780 460630 24808 699654
rect 41340 460698 41368 700402
rect 72988 700398 73016 703520
rect 89180 703474 89208 703520
rect 89364 703474 89392 703582
rect 89180 703446 89392 703474
rect 72976 700392 73028 700398
rect 72976 700334 73028 700340
rect 89640 460766 89668 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 154316 703582 154528 703610
rect 105464 700534 105492 703520
rect 137848 700670 137876 703520
rect 154132 703474 154160 703520
rect 154316 703474 154344 703582
rect 154132 703446 154344 703474
rect 137836 700664 137888 700670
rect 137836 700606 137888 700612
rect 105452 700528 105504 700534
rect 105452 700470 105504 700476
rect 106188 700528 106240 700534
rect 106188 700470 106240 700476
rect 106200 460834 106228 700470
rect 154500 460902 154528 703582
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 284036 703582 284248 703610
rect 170324 699718 170352 703520
rect 202800 700942 202828 703520
rect 218992 702434 219020 703520
rect 218992 702406 219388 702434
rect 202788 700936 202840 700942
rect 202788 700878 202840 700884
rect 170312 699712 170364 699718
rect 170312 699654 170364 699660
rect 171048 699712 171100 699718
rect 171048 699654 171100 699660
rect 154488 460896 154540 460902
rect 154488 460838 154540 460844
rect 106188 460828 106240 460834
rect 106188 460770 106240 460776
rect 89628 460760 89680 460766
rect 89628 460702 89680 460708
rect 41328 460692 41380 460698
rect 41328 460634 41380 460640
rect 24768 460624 24820 460630
rect 24768 460566 24820 460572
rect 3976 460216 4028 460222
rect 3976 460158 4028 460164
rect 171060 460154 171088 699654
rect 171048 460148 171100 460154
rect 171048 460090 171100 460096
rect 219360 460086 219388 702406
rect 235184 699718 235212 703520
rect 267660 700126 267688 703520
rect 283852 703474 283880 703520
rect 284036 703474 284064 703582
rect 283852 703446 284064 703474
rect 267648 700120 267700 700126
rect 267648 700062 267700 700068
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 235908 699712 235960 699718
rect 235908 699654 235960 699660
rect 219348 460080 219400 460086
rect 219348 460022 219400 460028
rect 235920 460018 235948 699654
rect 235908 460012 235960 460018
rect 235908 459954 235960 459960
rect 284220 459950 284248 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 300136 699718 300164 703520
rect 317328 701004 317380 701010
rect 317328 700946 317380 700952
rect 313188 700868 313240 700874
rect 313188 700810 313240 700816
rect 311808 700732 311860 700738
rect 311808 700674 311860 700680
rect 309048 700596 309100 700602
rect 309048 700538 309100 700544
rect 307668 700460 307720 700466
rect 307668 700402 307720 700408
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 300768 699712 300820 699718
rect 300768 699654 300820 699660
rect 299388 643136 299440 643142
rect 299388 643078 299440 643084
rect 298008 616888 298060 616894
rect 298008 616830 298060 616836
rect 295248 590708 295300 590714
rect 295248 590650 295300 590656
rect 293868 563100 293920 563106
rect 293868 563042 293920 563048
rect 289728 536852 289780 536858
rect 289728 536794 289780 536800
rect 288348 510672 288400 510678
rect 288348 510614 288400 510620
rect 285588 484424 285640 484430
rect 285588 484366 285640 484372
rect 284208 459944 284260 459950
rect 284208 459886 284260 459892
rect 281448 459740 281500 459746
rect 281448 459682 281500 459688
rect 272340 459604 272392 459610
rect 272340 459546 272392 459552
rect 255044 458856 255096 458862
rect 255044 458798 255096 458804
rect 228364 458584 228416 458590
rect 228364 458526 228416 458532
rect 222844 458448 222896 458454
rect 222844 458390 222896 458396
rect 3424 458244 3476 458250
rect 3424 458186 3476 458192
rect 3332 449880 3384 449886
rect 3332 449822 3384 449828
rect 3344 449585 3372 449822
rect 3330 449576 3386 449585
rect 3330 449511 3386 449520
rect 3436 423609 3464 458186
rect 4804 456816 4856 456822
rect 4804 456758 4856 456764
rect 3422 423600 3478 423609
rect 3422 423535 3478 423544
rect 3424 411256 3476 411262
rect 3424 411198 3476 411204
rect 3436 410553 3464 411198
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 3240 398812 3292 398818
rect 3240 398754 3292 398760
rect 3252 397497 3280 398754
rect 3238 397488 3294 397497
rect 3238 397423 3294 397432
rect 4816 371482 4844 456758
rect 222856 411262 222884 458390
rect 224224 457088 224276 457094
rect 224224 457030 224276 457036
rect 222844 411256 222896 411262
rect 222844 411198 222896 411204
rect 2780 371476 2832 371482
rect 2780 371418 2832 371424
rect 4804 371476 4856 371482
rect 4804 371418 4856 371424
rect 2792 371385 2820 371418
rect 2778 371376 2834 371385
rect 2778 371311 2834 371320
rect 224236 358766 224264 457030
rect 226984 457020 227036 457026
rect 226984 456962 227036 456968
rect 3332 358760 3384 358766
rect 3332 358702 3384 358708
rect 224224 358760 224276 358766
rect 224224 358702 224276 358708
rect 3344 358465 3372 358702
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3148 346384 3200 346390
rect 3148 346326 3200 346332
rect 3160 345409 3188 346326
rect 3146 345400 3202 345409
rect 3146 345335 3202 345344
rect 220084 336728 220136 336734
rect 220084 336670 220136 336676
rect 215944 336660 215996 336666
rect 215944 336602 215996 336608
rect 214564 336592 214616 336598
rect 214564 336534 214616 336540
rect 209044 336524 209096 336530
rect 209044 336466 209096 336472
rect 125508 336456 125560 336462
rect 43442 336424 43498 336433
rect 125508 336398 125560 336404
rect 43442 336359 43498 336368
rect 114468 336388 114520 336394
rect 25502 336288 25558 336297
rect 25502 336223 25558 336232
rect 18602 336152 18658 336161
rect 18602 336087 18658 336096
rect 7562 336016 7618 336025
rect 7562 335951 7618 335960
rect 3422 320104 3478 320113
rect 3422 320039 3478 320048
rect 3436 319297 3464 320039
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3330 293856 3386 293865
rect 3330 293791 3386 293800
rect 3344 293185 3372 293791
rect 3330 293176 3386 293185
rect 3330 293111 3386 293120
rect 3422 255232 3478 255241
rect 3422 255167 3478 255176
rect 3436 254153 3464 255167
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3422 202872 3478 202881
rect 3422 202807 3478 202816
rect 3436 201929 3464 202807
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 3422 164112 3478 164121
rect 3422 164047 3478 164056
rect 3436 162897 3464 164047
rect 3422 162888 3478 162897
rect 3422 162823 3478 162832
rect 3422 138000 3478 138009
rect 3422 137935 3478 137944
rect 3436 136785 3464 137935
rect 3422 136776 3478 136785
rect 3422 136711 3478 136720
rect 3422 111752 3478 111761
rect 3422 111687 3478 111696
rect 3436 110673 3464 111687
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 3422 85504 3478 85513
rect 3422 85439 3478 85448
rect 3436 84697 3464 85439
rect 3422 84688 3478 84697
rect 3422 84623 3478 84632
rect 3330 59256 3386 59265
rect 3330 59191 3386 59200
rect 3344 58585 3372 59191
rect 3330 58576 3386 58585
rect 3330 58511 3386 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3330 33144 3386 33153
rect 3330 33079 3386 33088
rect 3344 32473 3372 33079
rect 3330 32464 3386 32473
rect 3330 32399 3386 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4068 7608 4120 7614
rect 4068 7550 4120 7556
rect 2872 4956 2924 4962
rect 2872 4898 2924 4904
rect 1676 4888 1728 4894
rect 1676 4830 1728 4836
rect 572 4820 624 4826
rect 572 4762 624 4768
rect 584 480 612 4762
rect 1688 480 1716 4830
rect 2884 480 2912 4898
rect 4080 480 4108 7550
rect 7576 3874 7604 335951
rect 14464 327752 14516 327758
rect 14464 327694 14516 327700
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 5264 3868 5316 3874
rect 5264 3810 5316 3816
rect 7564 3868 7616 3874
rect 7564 3810 7616 3816
rect 5276 480 5304 3810
rect 6458 3360 6514 3369
rect 6458 3295 6514 3304
rect 6472 480 6500 3295
rect 7668 480 7696 4966
rect 8772 480 8800 8910
rect 12348 7676 12400 7682
rect 12348 7618 12400 7624
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 9956 2916 10008 2922
rect 9956 2858 10008 2864
rect 9968 480 9996 2858
rect 11164 480 11192 4082
rect 12360 480 12388 7618
rect 13544 3460 13596 3466
rect 13544 3402 13596 3408
rect 13556 480 13584 3402
rect 14476 2922 14504 327694
rect 17040 7744 17092 7750
rect 17040 7686 17092 7692
rect 15934 3632 15990 3641
rect 15934 3567 15990 3576
rect 14738 3496 14794 3505
rect 14738 3431 14794 3440
rect 14464 2916 14516 2922
rect 14464 2858 14516 2864
rect 14752 480 14780 3431
rect 15948 480 15976 3567
rect 17052 480 17080 7686
rect 18616 4146 18644 336087
rect 22744 334620 22796 334626
rect 22744 334562 22796 334568
rect 21824 7812 21876 7818
rect 21824 7754 21876 7760
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 20628 3664 20680 3670
rect 20628 3606 20680 3612
rect 18236 3596 18288 3602
rect 18236 3538 18288 3544
rect 18248 480 18276 3538
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 19444 480 19472 3334
rect 20640 480 20668 3606
rect 21836 480 21864 7754
rect 22756 3466 22784 334562
rect 24214 3768 24270 3777
rect 23020 3732 23072 3738
rect 24214 3703 24270 3712
rect 23020 3674 23072 3680
rect 22744 3460 22796 3466
rect 22744 3402 22796 3408
rect 23032 480 23060 3674
rect 24228 480 24256 3703
rect 25320 3460 25372 3466
rect 25320 3402 25372 3408
rect 25332 480 25360 3402
rect 25516 3398 25544 336223
rect 35164 336048 35216 336054
rect 35164 335990 35216 335996
rect 29644 334688 29696 334694
rect 29644 334630 29696 334636
rect 26516 7880 26568 7886
rect 26516 7822 26568 7828
rect 25504 3392 25556 3398
rect 25504 3334 25556 3340
rect 26528 480 26556 7822
rect 28908 3596 28960 3602
rect 28908 3538 28960 3544
rect 27712 3052 27764 3058
rect 27712 2994 27764 3000
rect 27724 480 27752 2994
rect 28920 480 28948 3538
rect 29656 3058 29684 334630
rect 33784 330540 33836 330546
rect 33784 330482 33836 330488
rect 32404 329180 32456 329186
rect 32404 329122 32456 329128
rect 30104 7948 30156 7954
rect 30104 7890 30156 7896
rect 29644 3052 29696 3058
rect 29644 2994 29696 3000
rect 30116 480 30144 7890
rect 32416 6914 32444 329122
rect 33600 9036 33652 9042
rect 33600 8978 33652 8984
rect 32324 6886 32444 6914
rect 32324 3534 32352 6886
rect 32312 3528 32364 3534
rect 32312 3470 32364 3476
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 31300 3392 31352 3398
rect 31300 3334 31352 3340
rect 31312 480 31340 3334
rect 32416 480 32444 3470
rect 33612 480 33640 8978
rect 33796 3398 33824 330482
rect 34796 4140 34848 4146
rect 34796 4082 34848 4088
rect 33784 3392 33836 3398
rect 33784 3334 33836 3340
rect 34808 480 34836 4082
rect 35176 3602 35204 335990
rect 39304 333260 39356 333266
rect 39304 333202 39356 333208
rect 36544 329112 36596 329118
rect 36544 329054 36596 329060
rect 36556 4146 36584 329054
rect 37188 9104 37240 9110
rect 37188 9046 37240 9052
rect 36544 4140 36596 4146
rect 36544 4082 36596 4088
rect 35992 3800 36044 3806
rect 35992 3742 36044 3748
rect 35164 3596 35216 3602
rect 35164 3538 35216 3544
rect 36004 480 36032 3742
rect 37200 480 37228 9046
rect 38384 3936 38436 3942
rect 38384 3878 38436 3884
rect 38396 480 38424 3878
rect 39316 3738 39344 333202
rect 41328 10328 41380 10334
rect 41328 10270 41380 10276
rect 39304 3732 39356 3738
rect 39304 3674 39356 3680
rect 39580 3664 39632 3670
rect 39580 3606 39632 3612
rect 39592 480 39620 3606
rect 41340 3602 41368 10270
rect 43076 4004 43128 4010
rect 43076 3946 43128 3952
rect 41880 3868 41932 3874
rect 41880 3810 41932 3816
rect 40684 3596 40736 3602
rect 40684 3538 40736 3544
rect 41328 3596 41380 3602
rect 41328 3538 41380 3544
rect 40696 480 40724 3538
rect 41892 480 41920 3810
rect 43088 480 43116 3946
rect 43456 3738 43484 336359
rect 114468 336330 114520 336336
rect 107568 336320 107620 336326
rect 107568 336262 107620 336268
rect 57244 336252 57296 336258
rect 57244 336194 57296 336200
rect 51724 336184 51776 336190
rect 51724 336126 51776 336132
rect 50344 336116 50396 336122
rect 50344 336058 50396 336064
rect 47584 329248 47636 329254
rect 47584 329190 47636 329196
rect 45468 10396 45520 10402
rect 45468 10338 45520 10344
rect 43444 3732 43496 3738
rect 43444 3674 43496 3680
rect 45376 3732 45428 3738
rect 45376 3674 45428 3680
rect 44272 3392 44324 3398
rect 44272 3334 44324 3340
rect 44284 480 44312 3334
rect 45388 1850 45416 3674
rect 45480 3398 45508 10338
rect 47596 3942 47624 329190
rect 49608 10464 49660 10470
rect 49608 10406 49660 10412
rect 47860 6180 47912 6186
rect 47860 6122 47912 6128
rect 47584 3936 47636 3942
rect 47584 3878 47636 3884
rect 45468 3392 45520 3398
rect 45468 3334 45520 3340
rect 46664 3392 46716 3398
rect 46664 3334 46716 3340
rect 45388 1822 45508 1850
rect 45480 480 45508 1822
rect 46676 480 46704 3334
rect 47872 480 47900 6122
rect 49620 3602 49648 10406
rect 50160 3936 50212 3942
rect 50160 3878 50212 3884
rect 48964 3596 49016 3602
rect 48964 3538 49016 3544
rect 49608 3596 49660 3602
rect 49608 3538 49660 3544
rect 48976 480 49004 3538
rect 50172 480 50200 3878
rect 50356 3806 50384 336058
rect 51356 6248 51408 6254
rect 51356 6190 51408 6196
rect 50344 3800 50396 3806
rect 50344 3742 50396 3748
rect 51368 480 51396 6190
rect 51736 4010 51764 336126
rect 54484 334756 54536 334762
rect 54484 334698 54536 334704
rect 53748 10532 53800 10538
rect 53748 10474 53800 10480
rect 51724 4004 51776 4010
rect 51724 3946 51776 3952
rect 53656 4004 53708 4010
rect 53656 3946 53708 3952
rect 52552 3596 52604 3602
rect 52552 3538 52604 3544
rect 52564 480 52592 3538
rect 53668 1986 53696 3946
rect 53760 3602 53788 10474
rect 54496 3874 54524 334698
rect 56508 10600 56560 10606
rect 56508 10542 56560 10548
rect 54944 6316 54996 6322
rect 54944 6258 54996 6264
rect 54484 3868 54536 3874
rect 54484 3810 54536 3816
rect 53748 3596 53800 3602
rect 53748 3538 53800 3544
rect 53668 1958 53788 1986
rect 53760 480 53788 1958
rect 54956 480 54984 6258
rect 56520 3398 56548 10542
rect 57256 4010 57284 336194
rect 86868 334892 86920 334898
rect 86868 334834 86920 334840
rect 84108 333328 84160 333334
rect 84108 333270 84160 333276
rect 68284 331900 68336 331906
rect 68284 331842 68336 331848
rect 61384 330608 61436 330614
rect 61384 330550 61436 330556
rect 58624 329316 58676 329322
rect 58624 329258 58676 329264
rect 58440 6384 58492 6390
rect 58440 6326 58492 6332
rect 57244 4004 57296 4010
rect 57244 3946 57296 3952
rect 56048 3392 56100 3398
rect 56048 3334 56100 3340
rect 56508 3392 56560 3398
rect 56508 3334 56560 3340
rect 56060 480 56088 3334
rect 57244 3188 57296 3194
rect 57244 3130 57296 3136
rect 57256 480 57284 3130
rect 58452 480 58480 6326
rect 58636 3738 58664 329258
rect 60648 10668 60700 10674
rect 60648 10610 60700 10616
rect 58624 3732 58676 3738
rect 58624 3674 58676 3680
rect 60660 3398 60688 10610
rect 60832 3732 60884 3738
rect 60832 3674 60884 3680
rect 59636 3392 59688 3398
rect 59636 3334 59688 3340
rect 60648 3392 60700 3398
rect 60648 3334 60700 3340
rect 59648 480 59676 3334
rect 60844 480 60872 3674
rect 61396 3194 61424 330550
rect 67548 10804 67600 10810
rect 67548 10746 67600 10752
rect 63224 10736 63276 10742
rect 63224 10678 63276 10684
rect 62028 6452 62080 6458
rect 62028 6394 62080 6400
rect 61384 3188 61436 3194
rect 61384 3130 61436 3136
rect 62040 480 62068 6394
rect 63236 480 63264 10678
rect 65524 6520 65576 6526
rect 65524 6462 65576 6468
rect 64328 3800 64380 3806
rect 64328 3742 64380 3748
rect 64340 480 64368 3742
rect 65536 480 65564 6462
rect 67560 3398 67588 10746
rect 68296 3942 68324 331842
rect 81348 330676 81400 330682
rect 81348 330618 81400 330624
rect 78588 11824 78640 11830
rect 78588 11766 78640 11772
rect 74448 11756 74500 11762
rect 74448 11698 74500 11704
rect 70308 10872 70360 10878
rect 70308 10814 70360 10820
rect 69112 6588 69164 6594
rect 69112 6530 69164 6536
rect 68284 3936 68336 3942
rect 68284 3878 68336 3884
rect 67916 3868 67968 3874
rect 67916 3810 67968 3816
rect 66720 3392 66772 3398
rect 66720 3334 66772 3340
rect 67548 3392 67600 3398
rect 67548 3334 67600 3340
rect 66732 480 66760 3334
rect 67928 480 67956 3810
rect 69124 480 69152 6530
rect 70320 480 70348 10814
rect 72608 8016 72660 8022
rect 72608 7958 72660 7964
rect 71504 3936 71556 3942
rect 71504 3878 71556 3884
rect 71516 480 71544 3878
rect 72620 480 72648 7958
rect 74460 3058 74488 11698
rect 76196 8084 76248 8090
rect 76196 8026 76248 8032
rect 75000 4004 75052 4010
rect 75000 3946 75052 3952
rect 73804 3052 73856 3058
rect 73804 2994 73856 3000
rect 74448 3052 74500 3058
rect 74448 2994 74500 3000
rect 73816 480 73844 2994
rect 75012 480 75040 3946
rect 76208 480 76236 8026
rect 78496 4140 78548 4146
rect 78496 4082 78548 4088
rect 77392 3392 77444 3398
rect 77392 3334 77444 3340
rect 77404 480 77432 3334
rect 78508 2122 78536 4082
rect 78600 3398 78628 11766
rect 79692 8152 79744 8158
rect 79692 8094 79744 8100
rect 78588 3392 78640 3398
rect 78588 3334 78640 3340
rect 78508 2094 78628 2122
rect 78600 480 78628 2094
rect 79704 480 79732 8094
rect 81360 3398 81388 330618
rect 82084 4072 82136 4078
rect 82084 4014 82136 4020
rect 80888 3392 80940 3398
rect 80888 3334 80940 3340
rect 81348 3392 81400 3398
rect 81348 3334 81400 3340
rect 80900 480 80928 3334
rect 82096 480 82124 4014
rect 84120 3398 84148 333270
rect 83280 3392 83332 3398
rect 83280 3334 83332 3340
rect 84108 3392 84160 3398
rect 84108 3334 84160 3340
rect 84476 3392 84528 3398
rect 84476 3334 84528 3340
rect 83292 480 83320 3334
rect 84488 480 84516 3334
rect 85672 3324 85724 3330
rect 85672 3266 85724 3272
rect 85684 480 85712 3266
rect 86880 480 86908 334834
rect 87604 334824 87656 334830
rect 87604 334766 87656 334772
rect 87616 3398 87644 334766
rect 104164 333532 104216 333538
rect 104164 333474 104216 333480
rect 93124 333464 93176 333470
rect 93124 333406 93176 333412
rect 88984 333396 89036 333402
rect 88984 333338 89036 333344
rect 88996 3398 89024 333338
rect 91008 10940 91060 10946
rect 91008 10882 91060 10888
rect 91020 3398 91048 10882
rect 93136 3398 93164 333406
rect 99288 332036 99340 332042
rect 99288 331978 99340 331984
rect 95148 331968 95200 331974
rect 95148 331910 95200 331916
rect 95056 11008 95108 11014
rect 95056 10950 95108 10956
rect 87604 3392 87656 3398
rect 87604 3334 87656 3340
rect 87972 3392 88024 3398
rect 87972 3334 88024 3340
rect 88984 3392 89036 3398
rect 88984 3334 89036 3340
rect 90364 3392 90416 3398
rect 90364 3334 90416 3340
rect 91008 3392 91060 3398
rect 91008 3334 91060 3340
rect 91560 3392 91612 3398
rect 91560 3334 91612 3340
rect 93124 3392 93176 3398
rect 93124 3334 93176 3340
rect 87984 480 88012 3334
rect 89168 3120 89220 3126
rect 89168 3062 89220 3068
rect 89180 480 89208 3062
rect 90376 480 90404 3334
rect 91572 480 91600 3334
rect 92756 3256 92808 3262
rect 92756 3198 92808 3204
rect 92768 480 92796 3198
rect 95068 3194 95096 10950
rect 93952 3188 94004 3194
rect 93952 3130 94004 3136
rect 95056 3188 95108 3194
rect 95056 3130 95108 3136
rect 93964 480 93992 3130
rect 95160 480 95188 331910
rect 97908 10260 97960 10266
rect 97908 10202 97960 10208
rect 97920 3330 97948 10202
rect 99300 3330 99328 331978
rect 102048 10192 102100 10198
rect 102048 10134 102100 10140
rect 102060 3330 102088 10134
rect 97448 3324 97500 3330
rect 97448 3266 97500 3272
rect 97908 3324 97960 3330
rect 97908 3266 97960 3272
rect 98644 3324 98696 3330
rect 98644 3266 98696 3272
rect 99288 3324 99340 3330
rect 99288 3266 99340 3272
rect 101036 3324 101088 3330
rect 101036 3266 101088 3272
rect 102048 3324 102100 3330
rect 102048 3266 102100 3272
rect 96252 3188 96304 3194
rect 96252 3130 96304 3136
rect 96264 480 96292 3130
rect 97460 480 97488 3266
rect 98656 480 98684 3266
rect 99840 2984 99892 2990
rect 99840 2926 99892 2932
rect 99852 480 99880 2926
rect 101048 480 101076 3266
rect 104176 3126 104204 333474
rect 106188 332104 106240 332110
rect 106188 332046 106240 332052
rect 104532 10124 104584 10130
rect 104532 10066 104584 10072
rect 102232 3120 102284 3126
rect 102232 3062 102284 3068
rect 104164 3120 104216 3126
rect 104164 3062 104216 3068
rect 102244 480 102272 3062
rect 103336 3052 103388 3058
rect 103336 2994 103388 3000
rect 103348 480 103376 2994
rect 104544 480 104572 10066
rect 106200 3126 106228 332046
rect 107580 3126 107608 336262
rect 113088 330812 113140 330818
rect 113088 330754 113140 330760
rect 111064 330744 111116 330750
rect 111064 330686 111116 330692
rect 108948 10056 109000 10062
rect 108948 9998 109000 10004
rect 108960 3126 108988 9998
rect 111076 3126 111104 330686
rect 111616 9988 111668 9994
rect 111616 9930 111668 9936
rect 105728 3120 105780 3126
rect 105728 3062 105780 3068
rect 106188 3120 106240 3126
rect 106188 3062 106240 3068
rect 106924 3120 106976 3126
rect 106924 3062 106976 3068
rect 107568 3120 107620 3126
rect 107568 3062 107620 3068
rect 108120 3120 108172 3126
rect 108120 3062 108172 3068
rect 108948 3120 109000 3126
rect 108948 3062 109000 3068
rect 109316 3120 109368 3126
rect 109316 3062 109368 3068
rect 111064 3120 111116 3126
rect 111064 3062 111116 3068
rect 105740 480 105768 3062
rect 106936 480 106964 3062
rect 108132 480 108160 3062
rect 109328 480 109356 3062
rect 110512 2984 110564 2990
rect 110512 2926 110564 2932
rect 110524 480 110552 2926
rect 111628 480 111656 9930
rect 113100 6914 113128 330754
rect 112824 6886 113128 6914
rect 112824 480 112852 6886
rect 114480 2922 114508 336330
rect 124128 332172 124180 332178
rect 124128 332114 124180 332120
rect 117228 330880 117280 330886
rect 117228 330822 117280 330828
rect 115848 9920 115900 9926
rect 115848 9862 115900 9868
rect 115860 2922 115888 9862
rect 117240 2922 117268 330822
rect 119988 329384 120040 329390
rect 119988 329326 120040 329332
rect 119804 9852 119856 9858
rect 119804 9794 119856 9800
rect 119816 2922 119844 9794
rect 120000 6914 120028 329326
rect 122748 9784 122800 9790
rect 122748 9726 122800 9732
rect 119908 6886 120028 6914
rect 114008 2916 114060 2922
rect 114008 2858 114060 2864
rect 114468 2916 114520 2922
rect 114468 2858 114520 2864
rect 115204 2916 115256 2922
rect 115204 2858 115256 2864
rect 115848 2916 115900 2922
rect 115848 2858 115900 2864
rect 116400 2916 116452 2922
rect 116400 2858 116452 2864
rect 117228 2916 117280 2922
rect 117228 2858 117280 2864
rect 118792 2916 118844 2922
rect 118792 2858 118844 2864
rect 119804 2916 119856 2922
rect 119804 2858 119856 2864
rect 114020 480 114048 2858
rect 115216 480 115244 2858
rect 116412 480 116440 2858
rect 117596 2848 117648 2854
rect 117596 2790 117648 2796
rect 117608 480 117636 2790
rect 118804 480 118832 2858
rect 119908 480 119936 6886
rect 121092 2848 121144 2854
rect 121092 2790 121144 2796
rect 121104 480 121132 2790
rect 122300 598 122512 626
rect 122300 480 122328 598
rect 122484 490 122512 598
rect 122760 490 122788 9726
rect 124140 6914 124168 332114
rect 125520 6914 125548 336398
rect 204904 335980 204956 335986
rect 204904 335922 204956 335928
rect 179328 335300 179380 335306
rect 179328 335242 179380 335248
rect 169668 335232 169720 335238
rect 169668 335174 169720 335180
rect 161388 335164 161440 335170
rect 161388 335106 161440 335112
rect 144828 335096 144880 335102
rect 144828 335038 144880 335044
rect 140688 334960 140740 334966
rect 140688 334902 140740 334908
rect 139308 15904 139360 15910
rect 139308 15846 139360 15852
rect 125876 13320 125928 13326
rect 125876 13262 125928 13268
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 122484 462 122788 490
rect 123496 6886 124168 6914
rect 125152 6886 125548 6914
rect 123496 480 123524 6886
rect 124692 598 124904 626
rect 124692 480 124720 598
rect 124876 490 124904 598
rect 125152 490 125180 6886
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 124876 462 125180 490
rect 125888 480 125916 13262
rect 128176 13116 128228 13122
rect 128176 13058 128228 13064
rect 126980 8900 127032 8906
rect 126980 8842 127032 8848
rect 126992 480 127020 8842
rect 128188 480 128216 13058
rect 135260 9240 135312 9246
rect 135260 9182 135312 9188
rect 131764 9172 131816 9178
rect 131764 9114 131816 9120
rect 130568 6656 130620 6662
rect 130568 6598 130620 6604
rect 129372 5092 129424 5098
rect 129372 5034 129424 5040
rect 129384 480 129412 5034
rect 130580 480 130608 6598
rect 131776 480 131804 9114
rect 134156 8220 134208 8226
rect 134156 8162 134208 8168
rect 132960 5160 133012 5166
rect 132960 5102 133012 5108
rect 132972 480 133000 5102
rect 134168 480 134196 8162
rect 135272 480 135300 9182
rect 137652 8288 137704 8294
rect 137652 8230 137704 8236
rect 136456 5296 136508 5302
rect 136456 5238 136508 5244
rect 136468 480 136496 5238
rect 137664 480 137692 8230
rect 138860 598 139072 626
rect 138860 480 138888 598
rect 139044 490 139072 598
rect 139320 490 139348 15846
rect 140700 6914 140728 334902
rect 143448 332240 143500 332246
rect 143448 332182 143500 332188
rect 141240 7540 141292 7546
rect 141240 7482 141292 7488
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 139044 462 139348 490
rect 140056 6886 140728 6914
rect 140056 480 140084 6886
rect 141252 480 141280 7482
rect 143460 6914 143488 332182
rect 144736 7472 144788 7478
rect 144736 7414 144788 7420
rect 142448 6886 143488 6914
rect 142448 480 142476 6886
rect 143540 4208 143592 4214
rect 143540 4150 143592 4156
rect 143552 480 143580 4150
rect 144748 480 144776 7414
rect 144840 4214 144868 335038
rect 147588 335028 147640 335034
rect 147588 334970 147640 334976
rect 146208 330948 146260 330954
rect 146208 330890 146260 330896
rect 146220 6914 146248 330890
rect 145944 6886 146248 6914
rect 144828 4208 144880 4214
rect 144828 4150 144880 4156
rect 145944 480 145972 6886
rect 147140 598 147352 626
rect 147140 480 147168 598
rect 147324 490 147352 598
rect 147600 490 147628 334970
rect 158628 333668 158680 333674
rect 158628 333610 158680 333616
rect 151728 333600 151780 333606
rect 151728 333542 151780 333548
rect 149980 13184 150032 13190
rect 149980 13126 150032 13132
rect 148324 7404 148376 7410
rect 148324 7346 148376 7352
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 147324 462 147628 490
rect 148336 480 148364 7346
rect 149532 598 149744 626
rect 149532 480 149560 598
rect 149716 490 149744 598
rect 149992 490 150020 13126
rect 151740 6914 151768 333542
rect 153108 331016 153160 331022
rect 153108 330958 153160 330964
rect 151820 7336 151872 7342
rect 151820 7278 151872 7284
rect 151096 6886 151768 6914
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 149716 462 150020 490
rect 150636 598 150848 626
rect 150636 480 150664 598
rect 150820 490 150848 598
rect 151096 490 151124 6886
rect 150594 -960 150706 480
rect 150820 462 151124 490
rect 151832 480 151860 7278
rect 153120 6914 153148 330958
rect 157248 18624 157300 18630
rect 157248 18566 157300 18572
rect 154212 11960 154264 11966
rect 154212 11902 154264 11908
rect 153028 6886 153148 6914
rect 153028 480 153056 6886
rect 154224 480 154252 11902
rect 155408 7268 155460 7274
rect 155408 7210 155460 7216
rect 155420 480 155448 7210
rect 157260 6914 157288 18566
rect 158640 6914 158668 333610
rect 161296 17264 161348 17270
rect 161296 17206 161348 17212
rect 161308 11694 161336 17206
rect 160100 11688 160152 11694
rect 160100 11630 160152 11636
rect 161296 11688 161348 11694
rect 161296 11630 161348 11636
rect 158904 7200 158956 7206
rect 158904 7142 158956 7148
rect 156616 6886 157288 6914
rect 158272 6886 158668 6914
rect 156616 480 156644 6886
rect 157812 598 158024 626
rect 157812 480 157840 598
rect 157996 490 158024 598
rect 158272 490 158300 6886
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 157996 462 158300 490
rect 158916 480 158944 7142
rect 160112 480 160140 11630
rect 161400 6914 161428 335106
rect 162768 333736 162820 333742
rect 162768 333678 162820 333684
rect 162780 6914 162808 333678
rect 164148 13252 164200 13258
rect 164148 13194 164200 13200
rect 161308 6886 161428 6914
rect 162504 6886 162808 6914
rect 161308 480 161336 6886
rect 162504 480 162532 6886
rect 163700 598 163912 626
rect 163700 480 163728 598
rect 163884 490 163912 598
rect 164160 490 164188 13194
rect 164884 12028 164936 12034
rect 164884 11970 164936 11976
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 163884 462 164188 490
rect 164896 480 164924 11970
rect 167644 11892 167696 11898
rect 167644 11834 167696 11840
rect 166080 6724 166132 6730
rect 166080 6666 166132 6672
rect 166092 480 166120 6666
rect 167196 598 167408 626
rect 167196 480 167224 598
rect 167380 490 167408 598
rect 167656 490 167684 11834
rect 169576 6792 169628 6798
rect 169576 6734 169628 6740
rect 168380 4208 168432 4214
rect 168380 4150 168432 4156
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 167380 462 167684 490
rect 168392 480 168420 4150
rect 169588 480 169616 6734
rect 169680 4214 169708 335174
rect 177948 333804 178000 333810
rect 177948 333746 178000 333752
rect 175188 332376 175240 332382
rect 175188 332318 175240 332324
rect 171048 332308 171100 332314
rect 171048 332250 171100 332256
rect 171060 6914 171088 332250
rect 175200 6914 175228 332318
rect 175924 12096 175976 12102
rect 175924 12038 175976 12044
rect 170784 6886 171088 6914
rect 174280 6886 175228 6914
rect 169668 4208 169720 4214
rect 169668 4150 169720 4156
rect 170784 480 170812 6886
rect 173164 6112 173216 6118
rect 173164 6054 173216 6060
rect 171968 4684 172020 4690
rect 171968 4626 172020 4632
rect 171980 480 172008 4626
rect 173176 480 173204 6054
rect 174280 480 174308 6886
rect 175476 598 175688 626
rect 175476 480 175504 598
rect 175660 490 175688 598
rect 175936 490 175964 12038
rect 177960 6914 177988 333746
rect 179340 6914 179368 335242
rect 197268 334552 197320 334558
rect 197268 334494 197320 334500
rect 188988 332512 189040 332518
rect 188988 332454 189040 332460
rect 182088 332444 182140 332450
rect 182088 332386 182140 332392
rect 182100 6914 182128 332386
rect 184940 13388 184992 13394
rect 184940 13330 184992 13336
rect 182548 12164 182600 12170
rect 182548 12106 182600 12112
rect 177868 6886 177988 6914
rect 179064 6886 179368 6914
rect 181456 6886 182128 6914
rect 176660 6044 176712 6050
rect 176660 5986 176712 5992
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 175660 462 175964 490
rect 176672 480 176700 5986
rect 177868 480 177896 6886
rect 179064 480 179092 6886
rect 180248 5976 180300 5982
rect 180248 5918 180300 5924
rect 180260 480 180288 5918
rect 181456 480 181484 6886
rect 182560 480 182588 12106
rect 183744 5908 183796 5914
rect 183744 5850 183796 5856
rect 183756 480 183784 5850
rect 184952 480 184980 13330
rect 187332 5840 187384 5846
rect 187332 5782 187384 5788
rect 186136 5500 186188 5506
rect 186136 5442 186188 5448
rect 186148 480 186176 5442
rect 187344 480 187372 5782
rect 188540 598 188752 626
rect 188540 480 188568 598
rect 188724 490 188752 598
rect 189000 490 189028 332454
rect 195612 9376 195664 9382
rect 195612 9318 195664 9324
rect 192024 9308 192076 9314
rect 192024 9250 192076 9256
rect 190828 5772 190880 5778
rect 190828 5714 190880 5720
rect 189724 5432 189776 5438
rect 189724 5374 189776 5380
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 188724 462 189028 490
rect 189736 480 189764 5374
rect 190840 480 190868 5714
rect 192036 480 192064 9250
rect 194416 5704 194468 5710
rect 194416 5646 194468 5652
rect 193220 4752 193272 4758
rect 193220 4694 193272 4700
rect 193232 480 193260 4694
rect 194428 480 194456 5646
rect 195624 480 195652 9318
rect 196820 598 197032 626
rect 196820 480 196848 598
rect 197004 490 197032 598
rect 197280 490 197308 334494
rect 202788 334484 202840 334490
rect 202788 334426 202840 334432
rect 198648 333872 198700 333878
rect 198648 333814 198700 333820
rect 198660 6914 198688 333814
rect 202696 9512 202748 9518
rect 202696 9454 202748 9460
rect 199108 9444 199160 9450
rect 199108 9386 199160 9392
rect 198384 6886 198688 6914
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197004 462 197308 490
rect 197924 598 198136 626
rect 197924 480 197952 598
rect 198108 490 198136 598
rect 198384 490 198412 6886
rect 197882 -960 197994 480
rect 198108 462 198412 490
rect 199120 480 199148 9386
rect 200304 4276 200356 4282
rect 200304 4218 200356 4224
rect 200316 480 200344 4218
rect 201500 4208 201552 4214
rect 201500 4150 201552 4156
rect 201512 480 201540 4150
rect 202708 480 202736 9454
rect 202800 4214 202828 334426
rect 204916 5302 204944 335922
rect 205548 333940 205600 333946
rect 205548 333882 205600 333888
rect 204904 5296 204956 5302
rect 204904 5238 204956 5244
rect 203892 5228 203944 5234
rect 203892 5170 203944 5176
rect 202788 4208 202840 4214
rect 202788 4150 202840 4156
rect 203904 480 203932 5170
rect 205100 598 205312 626
rect 205100 480 205128 598
rect 205284 490 205312 598
rect 205560 490 205588 333882
rect 209056 16574 209084 336466
rect 213184 335708 213236 335714
rect 213184 335650 213236 335656
rect 209688 333192 209740 333198
rect 209688 333134 209740 333140
rect 208964 16546 209084 16574
rect 206192 9580 206244 9586
rect 206192 9522 206244 9528
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 205284 462 205588 490
rect 206204 480 206232 9522
rect 207388 5296 207440 5302
rect 207388 5238 207440 5244
rect 207400 480 207428 5238
rect 208964 4282 208992 16546
rect 209700 6914 209728 333134
rect 212172 12232 212224 12238
rect 212172 12174 212224 12180
rect 209780 9648 209832 9654
rect 209780 9590 209832 9596
rect 209056 6886 209728 6914
rect 208952 4276 209004 4282
rect 208952 4218 209004 4224
rect 208596 598 208808 626
rect 208596 480 208624 598
rect 208780 490 208808 598
rect 209056 490 209084 6886
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 208780 462 209084 490
rect 209792 480 209820 9590
rect 210976 5364 211028 5370
rect 210976 5306 211028 5312
rect 210988 480 211016 5306
rect 212184 480 212212 12174
rect 213196 8906 213224 335650
rect 213184 8900 213236 8906
rect 213184 8842 213236 8848
rect 213368 8900 213420 8906
rect 213368 8842 213420 8848
rect 213380 480 213408 8842
rect 214576 6914 214604 336534
rect 214300 6886 214604 6914
rect 214300 5438 214328 6886
rect 215956 5506 215984 336602
rect 216588 334416 216640 334422
rect 216588 334358 216640 334364
rect 216600 6914 216628 334358
rect 219256 332580 219308 332586
rect 219256 332522 219308 332528
rect 216864 8832 216916 8838
rect 216864 8774 216916 8780
rect 216048 6886 216628 6914
rect 215944 5500 215996 5506
rect 215944 5442 215996 5448
rect 214288 5432 214340 5438
rect 214288 5374 214340 5380
rect 214472 5432 214524 5438
rect 214472 5374 214524 5380
rect 214484 480 214512 5374
rect 216048 3482 216076 6886
rect 215680 3454 216076 3482
rect 215680 480 215708 3454
rect 216876 480 216904 8774
rect 218060 5500 218112 5506
rect 218060 5442 218112 5448
rect 218072 480 218100 5442
rect 219268 480 219296 332522
rect 220096 4758 220124 336670
rect 224224 335912 224276 335918
rect 224224 335854 224276 335860
rect 222844 335776 222896 335782
rect 222844 335718 222896 335724
rect 220452 8764 220504 8770
rect 220452 8706 220504 8712
rect 220084 4752 220136 4758
rect 220084 4694 220136 4700
rect 220464 480 220492 8706
rect 221556 4752 221608 4758
rect 221556 4694 221608 4700
rect 221568 480 221596 4694
rect 222856 4690 222884 335718
rect 223488 334348 223540 334354
rect 223488 334290 223540 334296
rect 223500 6914 223528 334290
rect 224236 12170 224264 335854
rect 226996 45558 227024 456962
rect 228376 346390 228404 458526
rect 232596 458312 232648 458318
rect 232596 458254 232648 458260
rect 231124 457292 231176 457298
rect 231124 457234 231176 457240
rect 231136 398818 231164 457234
rect 231124 398812 231176 398818
rect 231124 398754 231176 398760
rect 228364 346384 228416 346390
rect 228364 346326 228416 346332
rect 228364 335640 228416 335646
rect 228364 335582 228416 335588
rect 227628 333124 227680 333130
rect 227628 333066 227680 333072
rect 226984 45552 227036 45558
rect 226984 45494 227036 45500
rect 224224 12164 224276 12170
rect 224224 12106 224276 12112
rect 223948 8696 224000 8702
rect 223948 8638 224000 8644
rect 223224 6886 223528 6914
rect 222844 4684 222896 4690
rect 222844 4626 222896 4632
rect 222764 598 222976 626
rect 222764 480 222792 598
rect 222948 490 222976 598
rect 223224 490 223252 6886
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 222948 462 223252 490
rect 223960 480 223988 8638
rect 227536 8628 227588 8634
rect 227536 8570 227588 8576
rect 225144 4684 225196 4690
rect 225144 4626 225196 4632
rect 225156 480 225184 4626
rect 226340 4208 226392 4214
rect 226340 4150 226392 4156
rect 226352 480 226380 4150
rect 227548 480 227576 8570
rect 227640 4214 227668 333066
rect 228376 12102 228404 335582
rect 231124 335572 231176 335578
rect 231124 335514 231176 335520
rect 228364 12096 228416 12102
rect 228364 12038 228416 12044
rect 231136 12034 231164 335514
rect 232504 335504 232556 335510
rect 232504 335446 232556 335452
rect 231124 12028 231176 12034
rect 231124 11970 231176 11976
rect 232516 11966 232544 335446
rect 232608 215286 232636 458254
rect 255056 457994 255084 458798
rect 270408 458516 270460 458522
rect 270408 458458 270460 458464
rect 254748 457966 255084 457994
rect 270420 457994 270448 458458
rect 272352 457994 272380 459546
rect 278688 458720 278740 458726
rect 278688 458662 278740 458668
rect 277032 458380 277084 458386
rect 277032 458322 277084 458328
rect 277044 457994 277072 458322
rect 278700 457994 278728 458662
rect 280068 458652 280120 458658
rect 280068 458594 280120 458600
rect 280080 457994 280108 458594
rect 270420 457966 270480 457994
rect 272044 457966 272380 457994
rect 276828 457966 277072 457994
rect 278392 457966 278728 457994
rect 279956 457966 280108 457994
rect 281460 457994 281488 459682
rect 285600 459678 285628 484366
rect 286968 470620 287020 470626
rect 286968 470562 287020 470568
rect 286980 460934 287008 470562
rect 288360 460934 288388 510614
rect 286704 460906 287008 460934
rect 288268 460906 288388 460934
rect 285036 459672 285088 459678
rect 285036 459614 285088 459620
rect 285588 459672 285640 459678
rect 285588 459614 285640 459620
rect 285048 457994 285076 459614
rect 286704 457994 286732 460906
rect 288268 457994 288296 460906
rect 289740 457994 289768 536794
rect 291108 524476 291160 524482
rect 291108 524418 291160 524424
rect 291120 457994 291148 524418
rect 293880 459746 293908 563042
rect 295260 459746 295288 590650
rect 296628 576904 296680 576910
rect 296628 576846 296680 576852
rect 296640 459746 296668 576846
rect 298020 460934 298048 616830
rect 299400 460934 299428 643078
rect 300676 630692 300728 630698
rect 300676 630634 300728 630640
rect 297744 460906 298048 460934
rect 299308 460906 299428 460934
rect 292948 459740 293000 459746
rect 292948 459682 293000 459688
rect 293868 459740 293920 459746
rect 293868 459682 293920 459688
rect 294512 459740 294564 459746
rect 294512 459682 294564 459688
rect 295248 459740 295300 459746
rect 295248 459682 295300 459688
rect 296076 459740 296128 459746
rect 296076 459682 296128 459688
rect 296628 459740 296680 459746
rect 296628 459682 296680 459688
rect 292960 457994 292988 459682
rect 294524 457994 294552 459682
rect 296088 457994 296116 459682
rect 297744 457994 297772 460906
rect 299308 457994 299336 460906
rect 300688 457994 300716 630634
rect 300780 459814 300808 699654
rect 304908 696992 304960 696998
rect 304908 696934 304960 696940
rect 302148 670744 302200 670750
rect 302148 670686 302200 670692
rect 300768 459808 300820 459814
rect 300768 459750 300820 459756
rect 302160 458266 302188 670686
rect 304920 459746 304948 696934
rect 306288 683188 306340 683194
rect 306288 683130 306340 683136
rect 306300 459746 306328 683130
rect 307680 459746 307708 700402
rect 309060 460934 309088 700538
rect 310428 700528 310480 700534
rect 310428 700470 310480 700476
rect 310440 460934 310468 700470
rect 308784 460906 309088 460934
rect 310348 460906 310468 460934
rect 303988 459740 304040 459746
rect 303988 459682 304040 459688
rect 304908 459740 304960 459746
rect 304908 459682 304960 459688
rect 305552 459740 305604 459746
rect 305552 459682 305604 459688
rect 306288 459740 306340 459746
rect 306288 459682 306340 459688
rect 307116 459740 307168 459746
rect 307116 459682 307168 459688
rect 307668 459740 307720 459746
rect 307668 459682 307720 459688
rect 281460 457966 281520 457994
rect 284740 457966 285076 457994
rect 286304 457966 286732 457994
rect 287868 457966 288296 457994
rect 289432 457966 289768 457994
rect 290996 457966 291148 457994
rect 292652 457966 292988 457994
rect 294216 457966 294552 457994
rect 295780 457966 296116 457994
rect 297344 457966 297772 457994
rect 298908 457966 299336 457994
rect 300472 457966 300716 457994
rect 302114 458238 302188 458266
rect 302114 457980 302142 458238
rect 304000 457994 304028 459682
rect 305564 457994 305592 459682
rect 307128 457994 307156 459682
rect 308784 457994 308812 460906
rect 310348 457994 310376 460906
rect 311820 457994 311848 700674
rect 313200 458266 313228 700810
rect 315948 700800 316000 700806
rect 315948 700742 316000 700748
rect 315960 459746 315988 700742
rect 317340 459746 317368 700946
rect 331312 700936 331364 700942
rect 331312 700878 331364 700884
rect 320088 700256 320140 700262
rect 320088 700198 320140 700204
rect 318708 700188 318760 700194
rect 318708 700130 318760 700136
rect 318720 459746 318748 700130
rect 320100 460934 320128 700198
rect 327080 700120 327132 700126
rect 327080 700062 327132 700068
rect 321468 700052 321520 700058
rect 321468 699994 321520 700000
rect 319824 460906 320128 460934
rect 315028 459740 315080 459746
rect 315028 459682 315080 459688
rect 315948 459740 316000 459746
rect 315948 459682 316000 459688
rect 316592 459740 316644 459746
rect 316592 459682 316644 459688
rect 317328 459740 317380 459746
rect 317328 459682 317380 459688
rect 318156 459740 318208 459746
rect 318156 459682 318208 459688
rect 318708 459740 318760 459746
rect 318708 459682 318760 459688
rect 303692 457966 304028 457994
rect 305256 457966 305592 457994
rect 306820 457966 307156 457994
rect 308384 457966 308812 457994
rect 309948 457966 310376 457994
rect 311604 457966 311848 457994
rect 313154 458238 313228 458266
rect 313154 457980 313182 458238
rect 315040 457994 315068 459682
rect 316604 457994 316632 459682
rect 318168 457994 318196 459682
rect 319824 457994 319852 460906
rect 321480 457994 321508 699994
rect 324228 699984 324280 699990
rect 324228 699926 324280 699932
rect 322848 699916 322900 699922
rect 322848 699858 322900 699864
rect 322860 457994 322888 699858
rect 324240 458266 324268 699926
rect 325700 459876 325752 459882
rect 325700 459818 325752 459824
rect 314732 457966 315068 457994
rect 316296 457966 316632 457994
rect 317860 457966 318196 457994
rect 319424 457966 319852 457994
rect 321080 457966 321508 457994
rect 322644 457966 322888 457994
rect 324194 458238 324268 458266
rect 324194 457980 324222 458238
rect 325712 457994 325740 459818
rect 327092 457994 327120 700062
rect 331324 480254 331352 700878
rect 332520 699922 332548 703520
rect 336740 700664 336792 700670
rect 336740 700606 336792 700612
rect 332508 699916 332560 699922
rect 332508 699858 332560 699864
rect 333244 618316 333296 618322
rect 333244 618258 333296 618264
rect 331324 480226 331720 480254
rect 330208 460012 330260 460018
rect 330208 459954 330260 459960
rect 328552 459944 328604 459950
rect 328552 459886 328604 459892
rect 328564 457994 328592 459886
rect 330220 457994 330248 459954
rect 331692 457994 331720 480226
rect 333256 460086 333284 618258
rect 334900 460148 334952 460154
rect 334900 460090 334952 460096
rect 333244 460080 333296 460086
rect 333244 460022 333296 460028
rect 333336 460012 333388 460018
rect 333336 459954 333388 459960
rect 333348 457994 333376 459954
rect 334912 457994 334940 460090
rect 336752 457994 336780 700606
rect 340880 700392 340932 700398
rect 340880 700334 340932 700340
rect 338764 565888 338816 565894
rect 338764 565830 338816 565836
rect 338776 460902 338804 565830
rect 340892 480254 340920 700334
rect 345020 700324 345072 700330
rect 345020 700266 345072 700272
rect 342904 514820 342956 514826
rect 342904 514762 342956 514768
rect 340892 480226 341196 480254
rect 338120 460896 338172 460902
rect 338120 460838 338172 460844
rect 338764 460896 338816 460902
rect 338764 460838 338816 460844
rect 338132 457994 338160 460838
rect 339684 460828 339736 460834
rect 339684 460770 339736 460776
rect 339696 457994 339724 460770
rect 341168 457994 341196 480226
rect 342916 460766 342944 514762
rect 345032 480254 345060 700266
rect 348804 699990 348832 703520
rect 364996 700058 365024 703520
rect 397472 700194 397500 703520
rect 413664 700262 413692 703520
rect 429856 701010 429884 703520
rect 429844 701004 429896 701010
rect 429844 700946 429896 700952
rect 462332 700874 462360 703520
rect 462320 700868 462372 700874
rect 462320 700810 462372 700816
rect 478524 700806 478552 703520
rect 478512 700800 478564 700806
rect 478512 700742 478564 700748
rect 494808 700738 494836 703520
rect 494796 700732 494848 700738
rect 494796 700674 494848 700680
rect 527192 700602 527220 703520
rect 527180 700596 527232 700602
rect 527180 700538 527232 700544
rect 543476 700534 543504 703520
rect 543464 700528 543516 700534
rect 543464 700470 543516 700476
rect 559668 700466 559696 703520
rect 559656 700460 559708 700466
rect 559656 700402 559708 700408
rect 413652 700256 413704 700262
rect 413652 700198 413704 700204
rect 397460 700188 397512 700194
rect 397460 700130 397512 700136
rect 364984 700052 365036 700058
rect 364984 699994 365036 700000
rect 348792 699984 348844 699990
rect 348792 699926 348844 699932
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 350540 656940 350592 656946
rect 350540 656882 350592 656888
rect 350552 480254 350580 656882
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 354680 605872 354732 605878
rect 354680 605814 354732 605820
rect 354692 480254 354720 605814
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 360200 553444 360252 553450
rect 360200 553386 360252 553392
rect 345032 480226 345888 480254
rect 350552 480226 350672 480254
rect 354692 480226 355364 480254
rect 342812 460760 342864 460766
rect 342812 460702 342864 460708
rect 342904 460760 342956 460766
rect 342904 460702 342956 460708
rect 342824 457994 342852 460702
rect 344376 460692 344428 460698
rect 344376 460634 344428 460640
rect 344388 457994 344416 460634
rect 345860 457994 345888 480226
rect 348516 462392 348568 462398
rect 348516 462334 348568 462340
rect 348528 460630 348556 462334
rect 347780 460624 347832 460630
rect 347780 460566 347832 460572
rect 348516 460624 348568 460630
rect 348516 460566 348568 460572
rect 347792 457994 347820 460566
rect 349160 460556 349212 460562
rect 349160 460498 349212 460504
rect 349172 457994 349200 460498
rect 350644 457994 350672 480226
rect 352288 460488 352340 460494
rect 352288 460430 352340 460436
rect 352300 457994 352328 460430
rect 353852 460420 353904 460426
rect 353852 460362 353904 460368
rect 353864 457994 353892 460362
rect 355336 457994 355364 480226
rect 358820 460352 358872 460358
rect 358820 460294 358872 460300
rect 356980 460080 357032 460086
rect 356980 460022 357032 460028
rect 356992 457994 357020 460022
rect 358832 457994 358860 460294
rect 360212 457994 360240 553386
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 364340 501016 364392 501022
rect 364340 500958 364392 500964
rect 364352 480254 364380 500958
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 364352 480226 364840 480254
rect 361764 460896 361816 460902
rect 361764 460838 361816 460844
rect 361776 457994 361804 460838
rect 363328 460284 363380 460290
rect 363328 460226 363380 460232
rect 363340 457994 363368 460226
rect 364812 457994 364840 480226
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 366456 460760 366508 460766
rect 366456 460702 366508 460708
rect 366468 457994 366496 460702
rect 371240 460624 371292 460630
rect 371240 460566 371292 460572
rect 368112 460216 368164 460222
rect 368112 460158 368164 460164
rect 368124 457994 368152 460158
rect 371252 457994 371280 460566
rect 556804 459672 556856 459678
rect 556804 459614 556856 459620
rect 555424 459604 555476 459610
rect 555424 459546 555476 459552
rect 418804 458720 418856 458726
rect 418804 458662 418856 458668
rect 379152 458584 379204 458590
rect 379152 458526 379204 458532
rect 375932 458448 375984 458454
rect 375932 458390 375984 458396
rect 373126 458244 373178 458250
rect 373126 458186 373178 458192
rect 325712 457966 325772 457994
rect 327092 457966 327336 457994
rect 328564 457966 328900 457994
rect 330220 457966 330556 457994
rect 331692 457966 332120 457994
rect 333348 457966 333684 457994
rect 334912 457966 335248 457994
rect 336752 457966 336812 457994
rect 338132 457966 338376 457994
rect 339696 457966 340032 457994
rect 341168 457966 341596 457994
rect 342824 457966 343160 457994
rect 344388 457966 344724 457994
rect 345860 457966 346288 457994
rect 347792 457966 347852 457994
rect 349172 457966 349508 457994
rect 350644 457966 351072 457994
rect 352300 457966 352636 457994
rect 353864 457966 354200 457994
rect 355336 457966 355764 457994
rect 356992 457966 357328 457994
rect 358832 457966 358984 457994
rect 360212 457966 360548 457994
rect 361776 457966 362112 457994
rect 363340 457966 363676 457994
rect 364812 457966 365240 457994
rect 366468 457966 366804 457994
rect 368124 457966 368460 457994
rect 371252 457966 371588 457994
rect 373138 457980 373166 458186
rect 375944 457994 375972 458390
rect 379164 457994 379192 458526
rect 391940 458312 391992 458318
rect 391940 458254 391992 458260
rect 391952 457994 391980 458254
rect 375944 457966 376280 457994
rect 379164 457966 379500 457994
rect 391952 457966 392104 457994
rect 238924 457434 239260 457450
rect 273700 457434 274036 457450
rect 275264 457434 275600 457450
rect 283176 457434 283512 457450
rect 233884 457428 233936 457434
rect 238924 457428 239272 457434
rect 238924 457422 239220 457428
rect 233884 457370 233936 457376
rect 273700 457428 274048 457434
rect 273700 457422 273996 457428
rect 239220 457370 239272 457376
rect 275264 457428 275612 457434
rect 275264 457422 275560 457428
rect 273996 457370 274048 457376
rect 283176 457428 283524 457434
rect 283176 457422 283472 457428
rect 275560 457370 275612 457376
rect 283472 457370 283524 457376
rect 233896 449886 233924 457370
rect 369860 457360 369912 457366
rect 237194 457328 237250 457337
rect 234632 457286 235796 457314
rect 233884 449880 233936 449886
rect 233884 449822 233936 449828
rect 233884 335844 233936 335850
rect 233884 335786 233936 335792
rect 232596 215280 232648 215286
rect 232596 215222 232648 215228
rect 233896 12238 233924 335786
rect 233976 335436 234028 335442
rect 233976 335378 234028 335384
rect 233988 13326 234016 335378
rect 233976 13320 234028 13326
rect 233976 13262 234028 13268
rect 233884 12232 233936 12238
rect 233884 12174 233936 12180
rect 232504 11960 232556 11966
rect 232504 11902 232556 11908
rect 231032 8560 231084 8566
rect 231032 8502 231084 8508
rect 229836 7132 229888 7138
rect 229836 7074 229888 7080
rect 228732 4616 228784 4622
rect 228732 4558 228784 4564
rect 227628 4208 227680 4214
rect 227628 4150 227680 4156
rect 228744 480 228772 4558
rect 229848 480 229876 7074
rect 231044 480 231072 8502
rect 233424 7064 233476 7070
rect 233424 7006 233476 7012
rect 232228 4548 232280 4554
rect 232228 4490 232280 4496
rect 232240 480 232268 4490
rect 233436 480 233464 7006
rect 234632 6866 234660 457286
rect 240782 457328 240838 457337
rect 237250 457286 237360 457314
rect 240488 457286 240782 457314
rect 237194 457263 237250 457272
rect 242346 457328 242402 457337
rect 242052 457286 242346 457314
rect 240782 457263 240838 457272
rect 243910 457328 243966 457337
rect 243616 457286 243910 457314
rect 242346 457263 242402 457272
rect 245474 457328 245530 457337
rect 245272 457286 245474 457314
rect 243910 457263 243966 457272
rect 246946 457328 247002 457337
rect 246836 457286 246946 457314
rect 245474 457263 245530 457272
rect 246946 457263 247002 457272
rect 248234 457328 248290 457337
rect 250258 457328 250314 457337
rect 248290 457286 248400 457314
rect 249964 457286 250258 457314
rect 248234 457263 248290 457272
rect 251822 457328 251878 457337
rect 251528 457286 251822 457314
rect 250258 457263 250314 457272
rect 253386 457328 253442 457337
rect 253092 457286 253386 457314
rect 251822 457263 251878 457272
rect 256514 457328 256570 457337
rect 256312 457286 256514 457314
rect 253386 457263 253442 457272
rect 256514 457263 256570 457272
rect 257526 457328 257582 457337
rect 259274 457328 259330 457337
rect 257582 457286 257876 457314
rect 257526 457263 257582 457272
rect 261298 457328 261354 457337
rect 259330 457286 259440 457314
rect 261004 457286 261298 457314
rect 259274 457263 259330 457272
rect 262862 457328 262918 457337
rect 262568 457286 262862 457314
rect 261298 457263 261354 457272
rect 264518 457328 264574 457337
rect 264224 457286 264518 457314
rect 262862 457263 262918 457272
rect 266082 457328 266138 457337
rect 265788 457286 266082 457314
rect 264518 457263 264574 457272
rect 267554 457328 267610 457337
rect 267352 457286 267554 457314
rect 266082 457263 266138 457272
rect 269026 457328 269082 457337
rect 268916 457286 269026 457314
rect 267554 457263 267610 457272
rect 374368 457360 374420 457366
rect 369912 457308 370024 457314
rect 369860 457302 370024 457308
rect 377588 457360 377640 457366
rect 374420 457308 374716 457314
rect 374368 457302 374716 457308
rect 380900 457360 380952 457366
rect 377640 457308 377936 457314
rect 377588 457302 377936 457308
rect 407580 457360 407632 457366
rect 382278 457328 382334 457337
rect 380952 457308 381064 457314
rect 380900 457302 381064 457308
rect 369872 457286 370024 457302
rect 374380 457286 374716 457302
rect 377600 457286 377936 457302
rect 380912 457286 381064 457302
rect 269026 457263 269082 457272
rect 384302 457328 384358 457337
rect 382334 457286 382628 457314
rect 384192 457286 384302 457314
rect 382278 457263 382334 457272
rect 384302 457263 384358 457272
rect 385406 457328 385462 457337
rect 387062 457328 387118 457337
rect 385462 457286 385756 457314
rect 385406 457263 385462 457272
rect 388626 457328 388682 457337
rect 387118 457286 387412 457314
rect 387062 457263 387118 457272
rect 390190 457328 390246 457337
rect 388682 457286 388976 457314
rect 388626 457263 388682 457272
rect 393502 457328 393558 457337
rect 390246 457286 390540 457314
rect 390190 457263 390246 457272
rect 394882 457328 394938 457337
rect 393558 457286 393668 457314
rect 393502 457263 393558 457272
rect 396538 457328 396594 457337
rect 394938 457286 395232 457314
rect 394882 457263 394938 457272
rect 398102 457328 398158 457337
rect 396594 457286 396888 457314
rect 396538 457263 396594 457272
rect 399666 457328 399722 457337
rect 398158 457286 398452 457314
rect 398102 457263 398158 457272
rect 401230 457328 401286 457337
rect 399722 457286 400016 457314
rect 399666 457263 399722 457272
rect 402978 457328 403034 457337
rect 401286 457286 401580 457314
rect 401230 457263 401286 457272
rect 404358 457328 404414 457337
rect 403034 457286 403144 457314
rect 402978 457263 403034 457272
rect 406014 457328 406070 457337
rect 404414 457286 404708 457314
rect 404358 457263 404414 457272
rect 406070 457286 406364 457314
rect 409142 457328 409198 457337
rect 407632 457308 407928 457314
rect 407580 457302 407928 457308
rect 407592 457286 407928 457302
rect 406014 457263 406070 457272
rect 410706 457328 410762 457337
rect 409198 457286 409492 457314
rect 409142 457263 409198 457272
rect 412270 457328 412326 457337
rect 410762 457286 411056 457314
rect 410706 457263 410762 457272
rect 412326 457286 412620 457314
rect 414184 457286 414980 457314
rect 412270 457263 412326 457272
rect 234908 338014 235152 338042
rect 235276 338014 235428 338042
rect 235552 338014 235796 338042
rect 234804 330472 234856 330478
rect 234804 330414 234856 330420
rect 234712 326324 234764 326330
rect 234712 326266 234764 326272
rect 234620 6860 234672 6866
rect 234620 6802 234672 6808
rect 234724 4962 234752 326266
rect 234712 4956 234764 4962
rect 234712 4898 234764 4904
rect 234816 4894 234844 330414
rect 234804 4888 234856 4894
rect 234804 4830 234856 4836
rect 234908 4826 234936 338014
rect 235276 330478 235304 338014
rect 235264 330472 235316 330478
rect 235264 330414 235316 330420
rect 235552 326330 235580 338014
rect 236150 337770 236178 338028
rect 236288 338014 236532 338042
rect 236656 338014 236900 338042
rect 237024 338014 237268 338042
rect 237484 338014 237636 338042
rect 237760 338014 238004 338042
rect 238128 338014 238372 338042
rect 238496 338014 238740 338042
rect 238864 338014 239108 338042
rect 239232 338014 239476 338042
rect 239600 338014 239844 338042
rect 240152 338014 240212 338042
rect 240336 338014 240580 338042
rect 240704 338014 240948 338042
rect 241072 338014 241316 338042
rect 236150 337742 236224 337770
rect 236092 330472 236144 330478
rect 236092 330414 236144 330420
rect 235540 326324 235592 326330
rect 235540 326266 235592 326272
rect 234988 8492 235040 8498
rect 234988 8434 235040 8440
rect 234896 4820 234948 4826
rect 234896 4762 234948 4768
rect 235000 3482 235028 8434
rect 236104 5030 236132 330414
rect 236196 7614 236224 337742
rect 236288 336025 236316 338014
rect 236274 336016 236330 336025
rect 236274 335951 236330 335960
rect 236656 316034 236684 338014
rect 237024 330478 237052 338014
rect 237012 330472 237064 330478
rect 237012 330414 237064 330420
rect 237380 330472 237432 330478
rect 237380 330414 237432 330420
rect 236288 316006 236684 316034
rect 236184 7608 236236 7614
rect 236184 7550 236236 7556
rect 236092 5024 236144 5030
rect 236092 4966 236144 4972
rect 235816 4820 235868 4826
rect 235816 4762 235868 4768
rect 234632 3454 235028 3482
rect 234632 480 234660 3454
rect 235828 480 235856 4762
rect 236288 3369 236316 316006
rect 237392 7682 237420 330414
rect 237484 8974 237512 338014
rect 237760 327758 237788 338014
rect 238128 336161 238156 338014
rect 238114 336152 238170 336161
rect 238114 336087 238170 336096
rect 238496 330478 238524 338014
rect 238864 334626 238892 338014
rect 239232 335354 239260 338014
rect 238956 335326 239260 335354
rect 238852 334620 238904 334626
rect 238852 334562 238904 334568
rect 238956 330528 238984 335326
rect 238864 330500 238984 330528
rect 238484 330472 238536 330478
rect 238484 330414 238536 330420
rect 237748 327752 237800 327758
rect 237748 327694 237800 327700
rect 237472 8968 237524 8974
rect 237472 8910 237524 8916
rect 238116 8968 238168 8974
rect 238116 8910 238168 8916
rect 237380 7676 237432 7682
rect 237380 7618 237432 7624
rect 237012 7608 237064 7614
rect 237012 7550 237064 7556
rect 236274 3360 236330 3369
rect 236274 3295 236330 3304
rect 237024 480 237052 7550
rect 238128 480 238156 8910
rect 238864 3505 238892 330500
rect 239600 316034 239628 338014
rect 238956 316006 239628 316034
rect 238956 3641 238984 316006
rect 240152 7750 240180 338014
rect 240336 329186 240364 338014
rect 240704 336297 240732 338014
rect 241072 336433 241100 338014
rect 241670 337770 241698 338028
rect 241808 338014 242052 338042
rect 242176 338014 242420 338042
rect 242544 338014 242788 338042
rect 243004 338014 243156 338042
rect 243280 338014 243524 338042
rect 243648 338014 243892 338042
rect 244016 338014 244260 338042
rect 244476 338014 244628 338042
rect 244752 338014 244996 338042
rect 245120 338014 245364 338042
rect 245672 338014 245732 338042
rect 245856 338014 246100 338042
rect 246224 338014 246468 338042
rect 246592 338014 246836 338042
rect 247112 338014 247264 338042
rect 241670 337742 241744 337770
rect 241058 336424 241114 336433
rect 241058 336359 241114 336368
rect 240690 336288 240746 336297
rect 240690 336223 240746 336232
rect 241612 330540 241664 330546
rect 241612 330482 241664 330488
rect 240324 329180 240376 329186
rect 240324 329122 240376 329128
rect 240140 7744 240192 7750
rect 240140 7686 240192 7692
rect 240508 7676 240560 7682
rect 240508 7618 240560 7624
rect 239312 4888 239364 4894
rect 239312 4830 239364 4836
rect 238942 3632 238998 3641
rect 238942 3567 238998 3576
rect 238850 3496 238906 3505
rect 238850 3431 238906 3440
rect 239324 480 239352 4830
rect 240520 480 240548 7618
rect 241624 3466 241652 330482
rect 241716 8514 241744 337742
rect 241808 333266 241836 338014
rect 241796 333260 241848 333266
rect 241796 333202 241848 333208
rect 242176 316034 242204 338014
rect 242544 330546 242572 338014
rect 242532 330540 242584 330546
rect 242532 330482 242584 330488
rect 241808 316006 242204 316034
rect 241808 16574 241836 316006
rect 241808 16546 241928 16574
rect 241716 8486 241836 8514
rect 241704 8424 241756 8430
rect 241704 8366 241756 8372
rect 241612 3460 241664 3466
rect 241612 3402 241664 3408
rect 241716 480 241744 8366
rect 241808 7818 241836 8486
rect 241796 7812 241848 7818
rect 241796 7754 241848 7760
rect 241900 3777 241928 16546
rect 243004 7886 243032 338014
rect 243280 334694 243308 338014
rect 243648 336054 243676 338014
rect 243636 336048 243688 336054
rect 243636 335990 243688 335996
rect 243268 334688 243320 334694
rect 243268 334630 243320 334636
rect 244016 316034 244044 338014
rect 244372 330540 244424 330546
rect 244372 330482 244424 330488
rect 243096 316006 244044 316034
rect 243096 7954 243124 316006
rect 244384 9042 244412 330482
rect 244476 330478 244504 338014
rect 244464 330472 244516 330478
rect 244464 330414 244516 330420
rect 244752 316034 244780 338014
rect 245120 330546 245148 338014
rect 245108 330540 245160 330546
rect 245108 330482 245160 330488
rect 245672 329118 245700 338014
rect 245856 336122 245884 338014
rect 245844 336116 245896 336122
rect 245844 336058 245896 336064
rect 245660 329112 245712 329118
rect 245660 329054 245712 329060
rect 246224 316034 246252 338014
rect 246592 329254 246620 338014
rect 247132 330540 247184 330546
rect 247132 330482 247184 330488
rect 246580 329248 246632 329254
rect 246580 329190 246632 329196
rect 244476 316006 244780 316034
rect 245948 316006 246252 316034
rect 244372 9036 244424 9042
rect 244372 8978 244424 8984
rect 243084 7948 243136 7954
rect 243084 7890 243136 7896
rect 242992 7880 243044 7886
rect 242992 7822 243044 7828
rect 244096 7744 244148 7750
rect 244096 7686 244148 7692
rect 242900 4956 242952 4962
rect 242900 4898 242952 4904
rect 241886 3768 241942 3777
rect 241886 3703 241942 3712
rect 242912 480 242940 4898
rect 244108 480 244136 7686
rect 244476 3534 244504 316006
rect 245948 9110 245976 316006
rect 247144 10334 247172 330482
rect 247132 10328 247184 10334
rect 247132 10270 247184 10276
rect 245936 9104 245988 9110
rect 245936 9046 245988 9052
rect 245200 9036 245252 9042
rect 245200 8978 245252 8984
rect 244464 3528 244516 3534
rect 244464 3470 244516 3476
rect 245212 480 245240 8978
rect 246396 5024 246448 5030
rect 246396 4966 246448 4972
rect 246408 480 246436 4966
rect 247236 3602 247264 338014
rect 247328 338014 247480 338042
rect 247604 338014 247848 338042
rect 247972 338014 248216 338042
rect 247328 330546 247356 338014
rect 247604 334762 247632 338014
rect 247972 336190 248000 338014
rect 248570 337770 248598 338028
rect 248708 338014 248952 338042
rect 249076 338014 249320 338042
rect 249444 338014 249688 338042
rect 249904 338014 250056 338042
rect 250180 338014 250424 338042
rect 250548 338014 250792 338042
rect 250916 338014 251160 338042
rect 251284 338014 251528 338042
rect 251652 338014 251896 338042
rect 252020 338014 252264 338042
rect 252572 338014 252632 338042
rect 252756 338014 253000 338042
rect 253124 338014 253368 338042
rect 253492 338014 253736 338042
rect 248570 337742 248644 337770
rect 247960 336184 248012 336190
rect 247960 336126 248012 336132
rect 247592 334756 247644 334762
rect 247592 334698 247644 334704
rect 247316 330540 247368 330546
rect 247316 330482 247368 330488
rect 248512 330540 248564 330546
rect 248512 330482 248564 330488
rect 247592 7812 247644 7818
rect 247592 7754 247644 7760
rect 247224 3596 247276 3602
rect 247224 3538 247276 3544
rect 247604 480 247632 7754
rect 248524 6186 248552 330482
rect 248616 10402 248644 337742
rect 248708 329322 248736 338014
rect 248696 329316 248748 329322
rect 248696 329258 248748 329264
rect 249076 316034 249104 338014
rect 249444 330546 249472 338014
rect 249432 330540 249484 330546
rect 249432 330482 249484 330488
rect 248708 316006 249104 316034
rect 248604 10396 248656 10402
rect 248604 10338 248656 10344
rect 248512 6180 248564 6186
rect 248512 6122 248564 6128
rect 248708 3670 248736 316006
rect 249904 10470 249932 338014
rect 250180 331906 250208 338014
rect 250168 331900 250220 331906
rect 250168 331842 250220 331848
rect 249984 330540 250036 330546
rect 249984 330482 250036 330488
rect 249996 10538 250024 330482
rect 250548 316034 250576 338014
rect 250916 330546 250944 338014
rect 251284 336258 251312 338014
rect 251272 336252 251324 336258
rect 251272 336194 251324 336200
rect 250904 330540 250956 330546
rect 250904 330482 250956 330488
rect 251272 330540 251324 330546
rect 251272 330482 251324 330488
rect 250088 316006 250576 316034
rect 249984 10532 250036 10538
rect 249984 10474 250036 10480
rect 249892 10464 249944 10470
rect 249892 10406 249944 10412
rect 248788 9104 248840 9110
rect 248788 9046 248840 9052
rect 248696 3664 248748 3670
rect 248696 3606 248748 3612
rect 248800 480 248828 9046
rect 250088 6254 250116 316006
rect 251088 11960 251140 11966
rect 251088 11902 251140 11908
rect 250076 6248 250128 6254
rect 250076 6190 250128 6196
rect 251100 3534 251128 11902
rect 251284 10606 251312 330482
rect 251652 316034 251680 338014
rect 252020 330546 252048 338014
rect 252572 330614 252600 338014
rect 252756 336682 252784 338014
rect 252664 336654 252784 336682
rect 252560 330608 252612 330614
rect 252560 330550 252612 330556
rect 252008 330540 252060 330546
rect 252008 330482 252060 330488
rect 251376 316006 251680 316034
rect 251272 10600 251324 10606
rect 251272 10542 251324 10548
rect 251180 7948 251232 7954
rect 251180 7890 251232 7896
rect 249984 3528 250036 3534
rect 249984 3470 250036 3476
rect 251088 3528 251140 3534
rect 251088 3470 251140 3476
rect 249996 480 250024 3470
rect 251192 480 251220 7890
rect 251376 6322 251404 316006
rect 252376 14476 252428 14482
rect 252376 14418 252428 14424
rect 251364 6316 251416 6322
rect 251364 6258 251416 6264
rect 252388 480 252416 14418
rect 252664 6390 252692 336654
rect 253124 335354 253152 338014
rect 252756 335326 253152 335354
rect 252756 10674 252784 335326
rect 253492 316034 253520 338014
rect 254090 337770 254118 338028
rect 254228 338014 254472 338042
rect 254596 338014 254840 338042
rect 254964 338014 255208 338042
rect 255516 338014 255576 338042
rect 255700 338014 255944 338042
rect 256068 338014 256312 338042
rect 256436 338014 256680 338042
rect 256804 338014 257048 338042
rect 257172 338014 257416 338042
rect 257540 338014 257784 338042
rect 258092 338014 258152 338042
rect 258276 338014 258520 338042
rect 258644 338014 258888 338042
rect 259012 338014 259164 338042
rect 254090 337742 254164 337770
rect 253940 330540 253992 330546
rect 253940 330482 253992 330488
rect 252848 316006 253520 316034
rect 252744 10668 252796 10674
rect 252744 10610 252796 10616
rect 252652 6384 252704 6390
rect 252652 6326 252704 6332
rect 252848 3738 252876 316006
rect 253848 10600 253900 10606
rect 253848 10542 253900 10548
rect 252836 3732 252888 3738
rect 252836 3674 252888 3680
rect 253492 598 253704 626
rect 253492 480 253520 598
rect 253676 490 253704 598
rect 253860 490 253888 10542
rect 253952 3806 253980 330482
rect 254032 330472 254084 330478
rect 254032 330414 254084 330420
rect 254044 6526 254072 330414
rect 254032 6520 254084 6526
rect 254032 6462 254084 6468
rect 254136 6458 254164 337742
rect 254228 10742 254256 338014
rect 254596 330546 254624 338014
rect 254584 330540 254636 330546
rect 254584 330482 254636 330488
rect 254964 330478 254992 338014
rect 255320 330540 255372 330546
rect 255320 330482 255372 330488
rect 254952 330472 255004 330478
rect 254952 330414 255004 330420
rect 254216 10736 254268 10742
rect 254216 10678 254268 10684
rect 254676 7880 254728 7886
rect 254676 7822 254728 7828
rect 254124 6452 254176 6458
rect 254124 6394 254176 6400
rect 253940 3800 253992 3806
rect 253940 3742 253992 3748
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 253676 462 253888 490
rect 254688 480 254716 7822
rect 255332 3874 255360 330482
rect 255412 330472 255464 330478
rect 255412 330414 255464 330420
rect 255424 6594 255452 330414
rect 255516 10810 255544 338014
rect 255700 330546 255728 338014
rect 255688 330540 255740 330546
rect 255688 330482 255740 330488
rect 256068 330478 256096 338014
rect 256056 330472 256108 330478
rect 256056 330414 256108 330420
rect 256436 316034 256464 338014
rect 256804 336682 256832 338014
rect 255608 316006 256464 316034
rect 256712 336654 256832 336682
rect 255608 10878 255636 316006
rect 255596 10872 255648 10878
rect 255596 10814 255648 10820
rect 255504 10804 255556 10810
rect 255504 10746 255556 10752
rect 256608 10328 256660 10334
rect 256608 10270 256660 10276
rect 255412 6588 255464 6594
rect 255412 6530 255464 6536
rect 255320 3868 255372 3874
rect 255320 3810 255372 3816
rect 256620 3534 256648 10270
rect 256712 3942 256740 336654
rect 257172 335354 257200 338014
rect 256804 335326 257200 335354
rect 256804 8022 256832 335326
rect 257540 316034 257568 338014
rect 256896 316006 257568 316034
rect 256896 11762 256924 316006
rect 256884 11756 256936 11762
rect 256884 11698 256936 11704
rect 256792 8016 256844 8022
rect 256792 7958 256844 7964
rect 257068 6180 257120 6186
rect 257068 6122 257120 6128
rect 256700 3936 256752 3942
rect 256700 3878 256752 3884
rect 255872 3528 255924 3534
rect 255872 3470 255924 3476
rect 256608 3528 256660 3534
rect 256608 3470 256660 3476
rect 255884 480 255912 3470
rect 257080 480 257108 6122
rect 258092 4010 258120 338014
rect 258172 330540 258224 330546
rect 258172 330482 258224 330488
rect 258184 4078 258212 330482
rect 258276 8242 258304 338014
rect 258644 316034 258672 338014
rect 259012 330546 259040 338014
rect 259518 337770 259546 338028
rect 259656 338014 259900 338042
rect 260024 338014 260268 338042
rect 260392 338014 260636 338042
rect 260944 338014 261004 338042
rect 261128 338014 261372 338042
rect 261496 338014 261740 338042
rect 261956 338014 262108 338042
rect 262324 338014 262476 338042
rect 262600 338014 262844 338042
rect 262968 338014 263212 338042
rect 263336 338014 263580 338042
rect 263704 338014 263948 338042
rect 264072 338014 264316 338042
rect 264440 338014 264684 338042
rect 259518 337742 259592 337770
rect 259460 336252 259512 336258
rect 259460 336194 259512 336200
rect 259472 334898 259500 336194
rect 259460 334892 259512 334898
rect 259460 334834 259512 334840
rect 259000 330540 259052 330546
rect 259000 330482 259052 330488
rect 258368 316006 258672 316034
rect 258368 11830 258396 316006
rect 258356 11824 258408 11830
rect 258356 11766 258408 11772
rect 258276 8214 258396 8242
rect 258368 8158 258396 8214
rect 259564 8158 259592 337742
rect 259656 330682 259684 338014
rect 259644 330676 259696 330682
rect 259644 330618 259696 330624
rect 260024 316034 260052 338014
rect 260392 333062 260420 338014
rect 260944 334830 260972 338014
rect 260932 334824 260984 334830
rect 260932 334766 260984 334772
rect 260380 333056 260432 333062
rect 260380 332998 260432 333004
rect 261128 316034 261156 338014
rect 261496 336258 261524 338014
rect 261484 336252 261536 336258
rect 261484 336194 261536 336200
rect 261956 333402 261984 338014
rect 261944 333396 261996 333402
rect 261944 333338 261996 333344
rect 259748 316006 260052 316034
rect 261036 316006 261156 316034
rect 258356 8152 258408 8158
rect 258356 8094 258408 8100
rect 259552 8152 259604 8158
rect 259552 8094 259604 8100
rect 258264 8084 258316 8090
rect 258264 8026 258316 8032
rect 258172 4072 258224 4078
rect 258172 4014 258224 4020
rect 258080 4004 258132 4010
rect 258080 3946 258132 3952
rect 258276 480 258304 8026
rect 259460 6316 259512 6322
rect 259460 6258 259512 6264
rect 259472 480 259500 6258
rect 259748 4146 259776 316006
rect 260656 10668 260708 10674
rect 260656 10610 260708 10616
rect 259736 4140 259788 4146
rect 259736 4082 259788 4088
rect 260668 480 260696 10610
rect 261036 3398 261064 316006
rect 261760 8084 261812 8090
rect 261760 8026 261812 8032
rect 261024 3392 261076 3398
rect 261024 3334 261076 3340
rect 261772 480 261800 8026
rect 262324 3330 262352 338014
rect 262600 335354 262628 338014
rect 262416 335326 262628 335354
rect 262416 10946 262444 335326
rect 262968 333470 262996 338014
rect 262956 333464 263008 333470
rect 262956 333406 263008 333412
rect 263336 316034 263364 338014
rect 263508 336048 263560 336054
rect 263508 335990 263560 335996
rect 262508 316006 263364 316034
rect 262404 10940 262456 10946
rect 262404 10882 262456 10888
rect 262312 3324 262364 3330
rect 262312 3266 262364 3272
rect 262508 3262 262536 316006
rect 263520 3534 263548 335990
rect 263704 11014 263732 338014
rect 264072 331974 264100 338014
rect 264060 331968 264112 331974
rect 264060 331910 264112 331916
rect 264440 316034 264468 338014
rect 265038 337770 265066 338028
rect 265176 338014 265420 338042
rect 265544 338014 265788 338042
rect 265912 338014 266156 338042
rect 266372 338014 266524 338042
rect 266648 338014 266892 338042
rect 267016 338014 267260 338042
rect 267384 338014 267628 338042
rect 267844 338014 267996 338042
rect 268120 338014 268364 338042
rect 268488 338014 268732 338042
rect 268856 338014 269100 338042
rect 269316 338014 269468 338042
rect 269592 338014 269836 338042
rect 269960 338014 270204 338042
rect 270572 338014 270724 338042
rect 265038 337742 265112 337770
rect 264888 336252 264940 336258
rect 264888 336194 264940 336200
rect 264900 332042 264928 336194
rect 264888 332036 264940 332042
rect 264888 331978 264940 331984
rect 263796 316006 264468 316034
rect 263692 11008 263744 11014
rect 263692 10950 263744 10956
rect 262956 3528 263008 3534
rect 262956 3470 263008 3476
rect 263508 3528 263560 3534
rect 263508 3470 263560 3476
rect 262496 3256 262548 3262
rect 262496 3198 262548 3204
rect 262968 480 262996 3470
rect 263796 3194 263824 316006
rect 264888 10396 264940 10402
rect 264888 10338 264940 10344
rect 264900 3534 264928 10338
rect 265084 10266 265112 337742
rect 265176 336258 265204 338014
rect 265164 336252 265216 336258
rect 265164 336194 265216 336200
rect 265164 330540 265216 330546
rect 265164 330482 265216 330488
rect 265072 10260 265124 10266
rect 265072 10202 265124 10208
rect 265176 10198 265204 330482
rect 265544 316034 265572 338014
rect 265912 330546 265940 338014
rect 266372 333538 266400 338014
rect 266360 333532 266412 333538
rect 266360 333474 266412 333480
rect 265900 330540 265952 330546
rect 265900 330482 265952 330488
rect 266452 330540 266504 330546
rect 266452 330482 266504 330488
rect 265268 316006 265572 316034
rect 265164 10192 265216 10198
rect 265164 10134 265216 10140
rect 264152 3528 264204 3534
rect 264152 3470 264204 3476
rect 264888 3528 264940 3534
rect 264888 3470 264940 3476
rect 263784 3188 263836 3194
rect 263784 3130 263836 3136
rect 264164 480 264192 3470
rect 265268 3126 265296 316006
rect 266464 10130 266492 330482
rect 266452 10124 266504 10130
rect 266452 10066 266504 10072
rect 265348 8152 265400 8158
rect 265348 8094 265400 8100
rect 265256 3120 265308 3126
rect 265256 3062 265308 3068
rect 265360 480 265388 8094
rect 266544 3528 266596 3534
rect 266544 3470 266596 3476
rect 266556 480 266584 3470
rect 266648 3058 266676 338014
rect 267016 330546 267044 338014
rect 267384 332110 267412 338014
rect 267844 336326 267872 338014
rect 267832 336320 267884 336326
rect 267832 336262 267884 336268
rect 267648 336184 267700 336190
rect 267648 336126 267700 336132
rect 267372 332104 267424 332110
rect 267372 332046 267424 332052
rect 267004 330540 267056 330546
rect 267004 330482 267056 330488
rect 267660 3534 267688 336126
rect 268120 335354 268148 338014
rect 267844 335326 268148 335354
rect 267844 10062 267872 335326
rect 268488 330750 268516 338014
rect 268476 330744 268528 330750
rect 268476 330686 268528 330692
rect 268856 316034 268884 338014
rect 269120 336252 269172 336258
rect 269120 336194 269172 336200
rect 269132 329390 269160 336194
rect 269120 329384 269172 329390
rect 269120 329326 269172 329332
rect 267936 316006 268884 316034
rect 267832 10056 267884 10062
rect 267832 9998 267884 10004
rect 267648 3528 267700 3534
rect 267648 3470 267700 3476
rect 267740 3528 267792 3534
rect 267740 3470 267792 3476
rect 266636 3052 266688 3058
rect 266636 2994 266688 3000
rect 267752 480 267780 3470
rect 267936 2990 267964 316006
rect 269028 10464 269080 10470
rect 269028 10406 269080 10412
rect 268844 6248 268896 6254
rect 268844 6190 268896 6196
rect 267924 2984 267976 2990
rect 267924 2926 267976 2932
rect 268856 480 268884 6190
rect 269040 3534 269068 10406
rect 269316 9994 269344 338014
rect 269592 330818 269620 338014
rect 269960 336394 269988 338014
rect 269948 336388 270000 336394
rect 269948 336330 270000 336336
rect 270408 336116 270460 336122
rect 270408 336058 270460 336064
rect 269580 330812 269632 330818
rect 269580 330754 269632 330760
rect 269304 9988 269356 9994
rect 269304 9930 269356 9936
rect 269028 3528 269080 3534
rect 269028 3470 269080 3476
rect 270052 598 270264 626
rect 270052 480 270080 598
rect 270236 490 270264 598
rect 270420 490 270448 336058
rect 270592 330540 270644 330546
rect 270592 330482 270644 330488
rect 270604 9858 270632 330482
rect 270696 9926 270724 338014
rect 270880 338014 270940 338042
rect 271064 338014 271216 338042
rect 271340 338014 271584 338042
rect 271892 338014 271952 338042
rect 272076 338014 272320 338042
rect 272444 338014 272688 338042
rect 272812 338014 273056 338042
rect 273272 338014 273424 338042
rect 273548 338014 273792 338042
rect 273916 338014 274160 338042
rect 274284 338014 274528 338042
rect 274652 338014 274896 338042
rect 275020 338014 275264 338042
rect 275388 338014 275632 338042
rect 275756 338014 276000 338042
rect 276216 338014 276368 338042
rect 276492 338014 276736 338042
rect 276860 338014 277104 338042
rect 270880 330886 270908 338014
rect 270868 330880 270920 330886
rect 270868 330822 270920 330828
rect 271064 316034 271092 338014
rect 271340 330546 271368 338014
rect 271788 336456 271840 336462
rect 271788 336398 271840 336404
rect 271800 332178 271828 336398
rect 271892 336258 271920 338014
rect 271880 336252 271932 336258
rect 271880 336194 271932 336200
rect 271788 332172 271840 332178
rect 271788 332114 271840 332120
rect 271328 330540 271380 330546
rect 271328 330482 271380 330488
rect 271972 330540 272024 330546
rect 271972 330482 272024 330488
rect 270788 316006 271092 316034
rect 270684 9920 270736 9926
rect 270684 9862 270736 9868
rect 270592 9852 270644 9858
rect 270592 9794 270644 9800
rect 270788 2922 270816 316006
rect 271788 10532 271840 10538
rect 271788 10474 271840 10480
rect 271800 3534 271828 10474
rect 271984 9790 272012 330482
rect 271972 9784 272024 9790
rect 271972 9726 272024 9732
rect 271236 3528 271288 3534
rect 271236 3470 271288 3476
rect 271788 3528 271840 3534
rect 271788 3470 271840 3476
rect 270776 2916 270828 2922
rect 270776 2858 270828 2864
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270236 462 270448 490
rect 271248 480 271276 3470
rect 272076 2854 272104 338014
rect 272444 330546 272472 338014
rect 272812 336462 272840 338014
rect 272800 336456 272852 336462
rect 272800 336398 272852 336404
rect 273272 336394 273300 338014
rect 273260 336388 273312 336394
rect 273260 336330 273312 336336
rect 273548 335442 273576 338014
rect 273916 335714 273944 338014
rect 273904 335708 273956 335714
rect 273904 335650 273956 335656
rect 273536 335436 273588 335442
rect 273536 335378 273588 335384
rect 272432 330540 272484 330546
rect 272432 330482 272484 330488
rect 274284 316034 274312 338014
rect 274548 336252 274600 336258
rect 274548 336194 274600 336200
rect 274456 335368 274508 335374
rect 274456 335310 274508 335316
rect 274468 332246 274496 335310
rect 274456 332240 274508 332246
rect 274456 332182 274508 332188
rect 273456 316006 274312 316034
rect 273456 13122 273484 316006
rect 273444 13116 273496 13122
rect 273444 13058 273496 13064
rect 274560 3534 274588 336194
rect 274652 5098 274680 338014
rect 275020 335354 275048 338014
rect 274836 335326 275048 335354
rect 274732 326392 274784 326398
rect 274732 326334 274784 326340
rect 274744 5166 274772 326334
rect 274836 6662 274864 335326
rect 275388 316034 275416 338014
rect 275756 326398 275784 338014
rect 276020 336456 276072 336462
rect 276020 336398 276072 336404
rect 276032 335102 276060 336398
rect 276020 335096 276072 335102
rect 276020 335038 276072 335044
rect 276216 326466 276244 338014
rect 276492 335354 276520 338014
rect 276860 335986 276888 338014
rect 277458 337770 277486 338028
rect 277596 338014 277840 338042
rect 277964 338014 278208 338042
rect 278332 338014 278576 338042
rect 278792 338014 278944 338042
rect 279068 338014 279312 338042
rect 279436 338014 279680 338042
rect 279804 338014 280048 338042
rect 280264 338014 280416 338042
rect 280540 338014 280784 338042
rect 280908 338014 281152 338042
rect 281460 338014 281520 338042
rect 281736 338014 281888 338042
rect 282012 338014 282256 338042
rect 282380 338014 282624 338042
rect 277458 337742 277532 337770
rect 277308 336388 277360 336394
rect 277308 336330 277360 336336
rect 276848 335980 276900 335986
rect 276848 335922 276900 335928
rect 276308 335326 276520 335354
rect 276204 326460 276256 326466
rect 276204 326402 276256 326408
rect 275744 326392 275796 326398
rect 275744 326334 275796 326340
rect 276204 326256 276256 326262
rect 276204 326198 276256 326204
rect 276112 321564 276164 321570
rect 276112 321506 276164 321512
rect 274928 316006 275416 316034
rect 274928 9178 274956 316006
rect 276124 9246 276152 321506
rect 276112 9240 276164 9246
rect 276112 9182 276164 9188
rect 274916 9172 274968 9178
rect 274916 9114 274968 9120
rect 276216 8226 276244 326198
rect 276308 321570 276336 335326
rect 276296 321564 276348 321570
rect 276296 321506 276348 321512
rect 276204 8220 276256 8226
rect 276204 8162 276256 8168
rect 274824 6656 274876 6662
rect 274824 6598 274876 6604
rect 274732 5160 274784 5166
rect 274732 5102 274784 5108
rect 274640 5092 274692 5098
rect 274640 5034 274692 5040
rect 274824 5092 274876 5098
rect 274824 5034 274876 5040
rect 273628 3528 273680 3534
rect 273628 3470 273680 3476
rect 274548 3528 274600 3534
rect 274548 3470 274600 3476
rect 272432 3460 272484 3466
rect 272432 3402 272484 3408
rect 272064 2848 272116 2854
rect 272064 2790 272116 2796
rect 272444 480 272472 3402
rect 273640 480 273668 3470
rect 274836 480 274864 5034
rect 277122 3360 277178 3369
rect 277122 3295 277178 3304
rect 276020 2916 276072 2922
rect 276020 2858 276072 2864
rect 276032 480 276060 2858
rect 277136 480 277164 3295
rect 277320 2922 277348 336330
rect 277504 326398 277532 337742
rect 277492 326392 277544 326398
rect 277492 326334 277544 326340
rect 277492 326256 277544 326262
rect 277492 326198 277544 326204
rect 277504 7546 277532 326198
rect 277596 15910 277624 338014
rect 277860 336456 277912 336462
rect 277860 336398 277912 336404
rect 277872 330954 277900 336398
rect 277964 334966 277992 338014
rect 277952 334960 278004 334966
rect 277952 334902 278004 334908
rect 277860 330948 277912 330954
rect 277860 330890 277912 330896
rect 277676 326392 277728 326398
rect 277676 326334 277728 326340
rect 277584 15904 277636 15910
rect 277584 15846 277636 15852
rect 277688 8294 277716 326334
rect 278332 326262 278360 338014
rect 278792 335374 278820 338014
rect 279068 336326 279096 338014
rect 279056 336320 279108 336326
rect 279056 336262 279108 336268
rect 278780 335368 278832 335374
rect 278780 335310 278832 335316
rect 278320 326256 278372 326262
rect 278320 326198 278372 326204
rect 279436 316034 279464 338014
rect 279804 336462 279832 338014
rect 279792 336456 279844 336462
rect 279792 336398 279844 336404
rect 280264 335034 280292 338014
rect 280252 335028 280304 335034
rect 280252 334970 280304 334976
rect 280252 326392 280304 326398
rect 280252 326334 280304 326340
rect 278976 316006 279464 316034
rect 277676 8288 277728 8294
rect 277676 8230 277728 8236
rect 277492 7540 277544 7546
rect 277492 7482 277544 7488
rect 278976 7478 279004 316006
rect 280264 13190 280292 326334
rect 280540 316034 280568 338014
rect 280908 326398 280936 338014
rect 281356 335980 281408 335986
rect 281356 335922 281408 335928
rect 281368 331214 281396 335922
rect 281460 333606 281488 338014
rect 281448 333600 281500 333606
rect 281448 333542 281500 333548
rect 281368 331186 281488 331214
rect 280896 326392 280948 326398
rect 280896 326334 280948 326340
rect 280356 316006 280568 316034
rect 280252 13184 280304 13190
rect 280252 13126 280304 13132
rect 278964 7472 279016 7478
rect 278964 7414 279016 7420
rect 280356 7410 280384 316006
rect 280344 7404 280396 7410
rect 280344 7346 280396 7352
rect 278320 5160 278372 5166
rect 278320 5102 278372 5108
rect 277308 2916 277360 2922
rect 277308 2858 277360 2864
rect 278332 480 278360 5102
rect 279516 3596 279568 3602
rect 279516 3538 279568 3544
rect 279528 480 279556 3538
rect 281460 3534 281488 331186
rect 281736 7342 281764 338014
rect 282012 331022 282040 338014
rect 282184 336320 282236 336326
rect 282184 336262 282236 336268
rect 282000 331016 282052 331022
rect 282000 330958 282052 330964
rect 282196 18630 282224 336262
rect 282380 335510 282408 338014
rect 282978 337770 283006 338028
rect 283116 338014 283268 338042
rect 283392 338014 283636 338042
rect 283760 338014 284004 338042
rect 282978 337742 283052 337770
rect 282644 336456 282696 336462
rect 282644 336398 282696 336404
rect 282368 335504 282420 335510
rect 282368 335446 282420 335452
rect 282656 333674 282684 336398
rect 282644 333668 282696 333674
rect 282644 333610 282696 333616
rect 282184 18624 282236 18630
rect 282184 18566 282236 18572
rect 281724 7336 281776 7342
rect 281724 7278 281776 7284
rect 283024 7274 283052 337742
rect 283116 336326 283144 338014
rect 283392 336462 283420 338014
rect 283380 336456 283432 336462
rect 283380 336398 283432 336404
rect 283104 336320 283156 336326
rect 283104 336262 283156 336268
rect 283760 316034 283788 338014
rect 284358 337770 284386 338028
rect 284496 338014 284740 338042
rect 284864 338014 285108 338042
rect 285232 338014 285476 338042
rect 285692 338014 285844 338042
rect 285968 338014 286212 338042
rect 286336 338014 286580 338042
rect 286704 338014 286948 338042
rect 287256 338014 287316 338042
rect 287440 338014 287684 338042
rect 287808 338014 288052 338042
rect 288176 338014 288420 338042
rect 288544 338014 288788 338042
rect 288912 338014 289156 338042
rect 289280 338014 289524 338042
rect 289832 338014 289892 338042
rect 290016 338014 290260 338042
rect 290384 338014 290628 338042
rect 290844 338014 290996 338042
rect 291212 338014 291364 338042
rect 291488 338014 291732 338042
rect 291856 338014 292100 338042
rect 292224 338014 292468 338042
rect 292684 338014 292836 338042
rect 292960 338014 293204 338042
rect 293328 338014 293572 338042
rect 293696 338014 293940 338042
rect 294064 338014 294308 338042
rect 294432 338014 294676 338042
rect 294800 338014 295044 338042
rect 295168 338014 295320 338042
rect 295444 338014 295688 338042
rect 295812 338014 296056 338042
rect 296180 338014 296424 338042
rect 296732 338014 296792 338042
rect 296916 338014 297160 338042
rect 297284 338014 297528 338042
rect 297652 338014 297896 338042
rect 298112 338014 298264 338042
rect 298388 338014 298632 338042
rect 298756 338014 299000 338042
rect 299124 338014 299368 338042
rect 299676 338014 299736 338042
rect 299860 338014 300104 338042
rect 300228 338014 300472 338042
rect 300596 338014 300840 338042
rect 301056 338014 301208 338042
rect 301332 338014 301576 338042
rect 301700 338014 301944 338042
rect 302312 338014 302556 338042
rect 284358 337742 284432 337770
rect 283116 316006 283788 316034
rect 283012 7268 283064 7274
rect 283012 7210 283064 7216
rect 283116 7206 283144 316006
rect 284404 17270 284432 337742
rect 284496 335170 284524 338014
rect 284484 335164 284536 335170
rect 284484 335106 284536 335112
rect 284864 333742 284892 338014
rect 284852 333736 284904 333742
rect 284852 333678 284904 333684
rect 285232 316034 285260 338014
rect 285692 335578 285720 338014
rect 285680 335572 285732 335578
rect 285680 335514 285732 335520
rect 285772 330540 285824 330546
rect 285772 330482 285824 330488
rect 284496 316006 285260 316034
rect 284392 17264 284444 17270
rect 284392 17206 284444 17212
rect 284496 13258 284524 316006
rect 284484 13252 284536 13258
rect 284484 13194 284536 13200
rect 285784 11898 285812 330482
rect 285968 316034 285996 338014
rect 286336 330546 286364 338014
rect 286416 335980 286468 335986
rect 286416 335922 286468 335928
rect 286324 330540 286376 330546
rect 286324 330482 286376 330488
rect 286428 316034 286456 335922
rect 286704 335238 286732 338014
rect 286692 335232 286744 335238
rect 286692 335174 286744 335180
rect 287152 330540 287204 330546
rect 287152 330482 287204 330488
rect 285876 316006 285996 316034
rect 286336 316006 286456 316034
rect 285772 11892 285824 11898
rect 285772 11834 285824 11840
rect 283104 7200 283156 7206
rect 283104 7142 283156 7148
rect 285876 6730 285904 316006
rect 286336 10674 286364 316006
rect 286324 10668 286376 10674
rect 286324 10610 286376 10616
rect 285864 6724 285916 6730
rect 285864 6666 285916 6672
rect 287164 6118 287192 330482
rect 287256 6798 287284 338014
rect 287440 332314 287468 338014
rect 287808 335782 287836 338014
rect 287796 335776 287848 335782
rect 287796 335718 287848 335724
rect 287428 332308 287480 332314
rect 287428 332250 287480 332256
rect 288176 330546 288204 338014
rect 288440 336728 288492 336734
rect 288440 336670 288492 336676
rect 288348 335708 288400 335714
rect 288348 335650 288400 335656
rect 288164 330540 288216 330546
rect 288164 330482 288216 330488
rect 287244 6792 287296 6798
rect 287244 6734 287296 6740
rect 287152 6112 287204 6118
rect 287152 6054 287204 6060
rect 281908 4480 281960 4486
rect 281908 4422 281960 4428
rect 280712 3528 280764 3534
rect 280712 3470 280764 3476
rect 281448 3528 281500 3534
rect 281448 3470 281500 3476
rect 280724 480 280752 3470
rect 281920 480 281948 4422
rect 285404 4412 285456 4418
rect 285404 4354 285456 4360
rect 284300 3596 284352 3602
rect 284300 3538 284352 3544
rect 283102 3496 283158 3505
rect 283102 3431 283158 3440
rect 283116 480 283144 3431
rect 284312 480 284340 3538
rect 285416 480 285444 4354
rect 286600 3664 286652 3670
rect 286600 3606 286652 3612
rect 286612 480 286640 3606
rect 288360 3398 288388 335650
rect 288452 333810 288480 336670
rect 288440 333804 288492 333810
rect 288440 333746 288492 333752
rect 288544 332382 288572 338014
rect 288912 335646 288940 338014
rect 289280 336682 289308 338014
rect 289832 336734 289860 338014
rect 289004 336654 289308 336682
rect 289820 336728 289872 336734
rect 289820 336670 289872 336676
rect 288900 335640 288952 335646
rect 288900 335582 288952 335588
rect 288532 332376 288584 332382
rect 288532 332318 288584 332324
rect 289004 316034 289032 336654
rect 289084 335776 289136 335782
rect 289084 335718 289136 335724
rect 288636 316006 289032 316034
rect 288636 6050 288664 316006
rect 289096 10606 289124 335718
rect 290016 335374 290044 338014
rect 290004 335368 290056 335374
rect 290004 335310 290056 335316
rect 290384 316034 290412 338014
rect 290844 332450 290872 338014
rect 291212 335918 291240 338014
rect 291200 335912 291252 335918
rect 291200 335854 291252 335860
rect 290832 332444 290884 332450
rect 290832 332386 290884 332392
rect 291292 330540 291344 330546
rect 291292 330482 291344 330488
rect 290016 316006 290412 316034
rect 289084 10600 289136 10606
rect 289084 10542 289136 10548
rect 288624 6044 288676 6050
rect 288624 5986 288676 5992
rect 290016 5982 290044 316006
rect 291304 13394 291332 330482
rect 291488 316034 291516 338014
rect 291568 336728 291620 336734
rect 291568 336670 291620 336676
rect 291580 332518 291608 336670
rect 291568 332512 291620 332518
rect 291568 332454 291620 332460
rect 291856 330546 291884 338014
rect 292224 336666 292252 338014
rect 292212 336660 292264 336666
rect 292212 336602 292264 336608
rect 292488 336660 292540 336666
rect 292488 336602 292540 336608
rect 291936 335912 291988 335918
rect 291936 335854 291988 335860
rect 291844 330540 291896 330546
rect 291844 330482 291896 330488
rect 291948 316034 291976 335854
rect 292500 334558 292528 336602
rect 292488 334552 292540 334558
rect 292488 334494 292540 334500
rect 291396 316006 291516 316034
rect 291856 316006 291976 316034
rect 291292 13388 291344 13394
rect 291292 13330 291344 13336
rect 290004 5976 290056 5982
rect 290004 5918 290056 5924
rect 291396 5914 291424 316006
rect 291856 11966 291884 316006
rect 291844 11960 291896 11966
rect 291844 11902 291896 11908
rect 291384 5908 291436 5914
rect 291384 5850 291436 5856
rect 292684 5846 292712 338014
rect 292960 336734 292988 338014
rect 292948 336728 293000 336734
rect 292948 336670 293000 336676
rect 293328 336598 293356 338014
rect 293316 336592 293368 336598
rect 293316 336534 293368 336540
rect 293696 316034 293724 338014
rect 292776 316006 293724 316034
rect 292672 5840 292724 5846
rect 292672 5782 292724 5788
rect 292776 5778 292804 316006
rect 294064 9314 294092 338014
rect 294432 336462 294460 338014
rect 294420 336456 294472 336462
rect 294420 336398 294472 336404
rect 294144 330540 294196 330546
rect 294144 330482 294196 330488
rect 294156 9382 294184 330482
rect 294800 316034 294828 338014
rect 295168 330546 295196 338014
rect 295444 336666 295472 338014
rect 295432 336660 295484 336666
rect 295432 336602 295484 336608
rect 295812 333878 295840 338014
rect 296180 336682 296208 338014
rect 295904 336654 296208 336682
rect 296536 336660 296588 336666
rect 295800 333872 295852 333878
rect 295800 333814 295852 333820
rect 295156 330540 295208 330546
rect 295156 330482 295208 330488
rect 295904 316034 295932 336654
rect 296536 336602 296588 336608
rect 295984 335708 296036 335714
rect 295984 335650 296036 335656
rect 294248 316006 294828 316034
rect 295536 316006 295932 316034
rect 294144 9376 294196 9382
rect 294144 9318 294196 9324
rect 294052 9308 294104 9314
rect 294052 9250 294104 9256
rect 292764 5772 292816 5778
rect 292764 5714 292816 5720
rect 294248 5710 294276 316006
rect 295536 9450 295564 316006
rect 295524 9444 295576 9450
rect 295524 9386 295576 9392
rect 295996 6322 296024 335650
rect 296444 335640 296496 335646
rect 296444 335582 296496 335588
rect 296456 333946 296484 335582
rect 296548 334490 296576 336602
rect 296628 336592 296680 336598
rect 296628 336534 296680 336540
rect 296536 334484 296588 334490
rect 296536 334426 296588 334432
rect 296444 333940 296496 333946
rect 296444 333882 296496 333888
rect 295984 6316 296036 6322
rect 295984 6258 296036 6264
rect 294236 5704 294288 5710
rect 294236 5646 294288 5652
rect 288992 4344 289044 4350
rect 288992 4286 289044 4292
rect 287796 3392 287848 3398
rect 287796 3334 287848 3340
rect 288348 3392 288400 3398
rect 288348 3334 288400 3340
rect 287808 480 287836 3334
rect 289004 480 289032 4286
rect 292580 4276 292632 4282
rect 292580 4218 292632 4224
rect 291384 3732 291436 3738
rect 291384 3674 291436 3680
rect 290186 3632 290242 3641
rect 290186 3567 290242 3576
rect 290200 480 290228 3567
rect 291396 480 291424 3674
rect 292592 480 292620 4218
rect 293684 3800 293736 3806
rect 293684 3742 293736 3748
rect 294878 3768 294934 3777
rect 293696 480 293724 3742
rect 294878 3703 294934 3712
rect 294892 480 294920 3703
rect 296640 3058 296668 336534
rect 296732 336530 296760 338014
rect 296916 336666 296944 338014
rect 296904 336660 296956 336666
rect 296904 336602 296956 336608
rect 296720 336524 296772 336530
rect 296720 336466 296772 336472
rect 297284 335354 297312 338014
rect 296824 335326 297312 335354
rect 296824 9518 296852 335326
rect 297652 316034 297680 338014
rect 298112 335646 298140 338014
rect 298100 335640 298152 335646
rect 298100 335582 298152 335588
rect 298388 335354 298416 338014
rect 296916 316006 297680 316034
rect 298204 335326 298416 335354
rect 296812 9512 296864 9518
rect 296812 9454 296864 9460
rect 296916 5234 296944 316006
rect 298204 9586 298232 335326
rect 298756 316034 298784 338014
rect 299124 333198 299152 338014
rect 299388 336524 299440 336530
rect 299388 336466 299440 336472
rect 299112 333192 299164 333198
rect 299112 333134 299164 333140
rect 298296 316006 298784 316034
rect 298192 9580 298244 9586
rect 298192 9522 298244 9528
rect 298296 5302 298324 316006
rect 298284 5296 298336 5302
rect 298284 5238 298336 5244
rect 296904 5228 296956 5234
rect 296904 5170 296956 5176
rect 297272 3868 297324 3874
rect 297272 3810 297324 3816
rect 296076 3052 296128 3058
rect 296076 2994 296128 3000
rect 296628 3052 296680 3058
rect 296628 2994 296680 3000
rect 296088 480 296116 2994
rect 297284 480 297312 3810
rect 299400 3398 299428 336466
rect 299572 330540 299624 330546
rect 299572 330482 299624 330488
rect 299584 8906 299612 330482
rect 299676 9654 299704 338014
rect 299860 316034 299888 338014
rect 300228 335850 300256 338014
rect 300492 336728 300544 336734
rect 300492 336670 300544 336676
rect 300216 335844 300268 335850
rect 300216 335786 300268 335792
rect 300504 334422 300532 336670
rect 300492 334416 300544 334422
rect 300492 334358 300544 334364
rect 300596 330546 300624 338014
rect 300768 336660 300820 336666
rect 300768 336602 300820 336608
rect 300584 330540 300636 330546
rect 300584 330482 300636 330488
rect 299768 316006 299888 316034
rect 299664 9648 299716 9654
rect 299664 9590 299716 9596
rect 299572 8900 299624 8906
rect 299572 8842 299624 8848
rect 299664 6384 299716 6390
rect 299664 6326 299716 6332
rect 298468 3392 298520 3398
rect 298468 3334 298520 3340
rect 299388 3392 299440 3398
rect 299388 3334 299440 3340
rect 298480 480 298508 3334
rect 299676 480 299704 6326
rect 299768 5370 299796 316006
rect 299756 5364 299808 5370
rect 299756 5306 299808 5312
rect 300780 480 300808 336602
rect 300952 330540 301004 330546
rect 300952 330482 301004 330488
rect 300964 8838 300992 330482
rect 300952 8832 301004 8838
rect 300952 8774 301004 8780
rect 301056 5438 301084 338014
rect 301332 336734 301360 338014
rect 301320 336728 301372 336734
rect 301320 336670 301372 336676
rect 301700 330546 301728 338014
rect 301688 330540 301740 330546
rect 301688 330482 301740 330488
rect 302528 326466 302556 338014
rect 302620 338014 302680 338042
rect 302804 338014 303048 338042
rect 303172 338014 303416 338042
rect 303632 338014 303784 338042
rect 303908 338014 304152 338042
rect 304276 338014 304520 338042
rect 304644 338014 304888 338042
rect 305196 338014 305256 338042
rect 305380 338014 305624 338042
rect 305748 338014 305992 338042
rect 306116 338014 306360 338042
rect 306484 338014 306728 338042
rect 306852 338014 307096 338042
rect 307220 338014 307372 338042
rect 307496 338014 307740 338042
rect 307864 338014 308108 338042
rect 308232 338014 308476 338042
rect 308600 338014 308844 338042
rect 309212 338014 309364 338042
rect 302620 332586 302648 338014
rect 302804 335354 302832 338014
rect 302712 335326 302832 335354
rect 302608 332580 302660 332586
rect 302608 332522 302660 332528
rect 302712 331214 302740 335326
rect 302620 331186 302740 331214
rect 302516 326460 302568 326466
rect 302516 326402 302568 326408
rect 302332 326392 302384 326398
rect 302332 326334 302384 326340
rect 301044 5432 301096 5438
rect 301044 5374 301096 5380
rect 302344 4758 302372 326334
rect 302620 323762 302648 331186
rect 303172 326398 303200 338014
rect 303632 334354 303660 338014
rect 303908 335354 303936 338014
rect 303724 335326 303936 335354
rect 303620 334348 303672 334354
rect 303620 334290 303672 334296
rect 303160 326392 303212 326398
rect 303160 326334 303212 326340
rect 302436 323734 302648 323762
rect 302436 8770 302464 323734
rect 302516 323604 302568 323610
rect 302516 323546 302568 323552
rect 302424 8764 302476 8770
rect 302424 8706 302476 8712
rect 302528 5506 302556 323546
rect 303724 8702 303752 335326
rect 304276 316034 304304 338014
rect 304644 333130 304672 338014
rect 304908 336728 304960 336734
rect 304908 336670 304960 336676
rect 304632 333124 304684 333130
rect 304632 333066 304684 333072
rect 303816 316006 304304 316034
rect 303712 8696 303764 8702
rect 303712 8638 303764 8644
rect 303160 6316 303212 6322
rect 303160 6258 303212 6264
rect 302516 5500 302568 5506
rect 302516 5442 302568 5448
rect 302332 4752 302384 4758
rect 302332 4694 302384 4700
rect 301964 3936 302016 3942
rect 301964 3878 302016 3884
rect 301976 480 302004 3878
rect 303172 480 303200 6258
rect 303816 4690 303844 316006
rect 303804 4684 303856 4690
rect 303804 4626 303856 4632
rect 304920 3398 304948 336670
rect 305000 326392 305052 326398
rect 305000 326334 305052 326340
rect 305196 326346 305224 338014
rect 305380 326398 305408 338014
rect 305368 326392 305420 326398
rect 305012 4622 305040 326334
rect 305196 326318 305316 326346
rect 305368 326334 305420 326340
rect 305092 326256 305144 326262
rect 305092 326198 305144 326204
rect 305104 7138 305132 326198
rect 305184 326188 305236 326194
rect 305184 326130 305236 326136
rect 305196 8566 305224 326130
rect 305288 8634 305316 326318
rect 305748 326262 305776 338014
rect 305736 326256 305788 326262
rect 305736 326198 305788 326204
rect 306116 326194 306144 338014
rect 306380 326392 306432 326398
rect 306380 326334 306432 326340
rect 306104 326188 306156 326194
rect 306104 326130 306156 326136
rect 305276 8628 305328 8634
rect 305276 8570 305328 8576
rect 305184 8560 305236 8566
rect 305184 8502 305236 8508
rect 305092 7132 305144 7138
rect 305092 7074 305144 7080
rect 306392 4826 306420 326334
rect 306380 4820 306432 4826
rect 306380 4762 306432 4768
rect 305000 4616 305052 4622
rect 305000 4558 305052 4564
rect 306484 4554 306512 338014
rect 306852 335354 306880 338014
rect 306576 335326 306880 335354
rect 306576 7070 306604 335326
rect 307220 316034 307248 338014
rect 307496 326398 307524 338014
rect 307484 326392 307536 326398
rect 307484 326334 307536 326340
rect 307760 326392 307812 326398
rect 307760 326334 307812 326340
rect 306668 316006 307248 316034
rect 306668 8498 306696 316006
rect 306656 8492 306708 8498
rect 306656 8434 306708 8440
rect 306564 7064 306616 7070
rect 306564 7006 306616 7012
rect 307772 4894 307800 326334
rect 307864 7614 307892 338014
rect 308232 316034 308260 338014
rect 308600 326398 308628 338014
rect 309232 326460 309284 326466
rect 309232 326402 309284 326408
rect 308588 326392 308640 326398
rect 308588 326334 308640 326340
rect 309140 326392 309192 326398
rect 309140 326334 309192 326340
rect 307956 316006 308260 316034
rect 307956 8974 307984 316006
rect 307944 8968 307996 8974
rect 307944 8910 307996 8916
rect 307852 7608 307904 7614
rect 307852 7550 307904 7556
rect 309152 4962 309180 326334
rect 309244 7750 309272 326402
rect 309232 7744 309284 7750
rect 309232 7686 309284 7692
rect 309336 7682 309364 338014
rect 309428 338014 309580 338042
rect 309704 338014 309948 338042
rect 310072 338014 310316 338042
rect 309428 8430 309456 338014
rect 309704 326398 309732 338014
rect 310072 326466 310100 338014
rect 310670 337770 310698 338028
rect 310808 338014 311052 338042
rect 311176 338014 311420 338042
rect 311544 338014 311788 338042
rect 311912 338014 312156 338042
rect 312280 338014 312524 338042
rect 312648 338014 312892 338042
rect 313016 338014 313260 338042
rect 313384 338014 313628 338042
rect 313752 338014 313996 338042
rect 314120 338014 314364 338042
rect 314732 338014 314884 338042
rect 310670 337742 310744 337770
rect 310520 335708 310572 335714
rect 310520 335650 310572 335656
rect 310060 326460 310112 326466
rect 310060 326402 310112 326408
rect 309692 326392 309744 326398
rect 309692 326334 309744 326340
rect 309416 8424 309468 8430
rect 309416 8366 309468 8372
rect 309324 7676 309376 7682
rect 309324 7618 309376 7624
rect 310532 5030 310560 335650
rect 310612 326392 310664 326398
rect 310612 326334 310664 326340
rect 310624 7818 310652 326334
rect 310716 9042 310744 337742
rect 310808 335714 310836 338014
rect 310796 335708 310848 335714
rect 310796 335650 310848 335656
rect 311176 326398 311204 338014
rect 311164 326392 311216 326398
rect 311164 326334 311216 326340
rect 311544 316034 311572 338014
rect 311912 335918 311940 338014
rect 311900 335912 311952 335918
rect 311900 335854 311952 335860
rect 311992 330540 312044 330546
rect 311992 330482 312044 330488
rect 310808 316006 311572 316034
rect 310808 9110 310836 316006
rect 312004 14482 312032 330482
rect 312280 316034 312308 338014
rect 312648 330546 312676 338014
rect 313016 335782 313044 338014
rect 313004 335776 313056 335782
rect 313004 335718 313056 335724
rect 312636 330540 312688 330546
rect 312636 330482 312688 330488
rect 313280 330540 313332 330546
rect 313280 330482 313332 330488
rect 312096 316006 312308 316034
rect 311992 14476 312044 14482
rect 311992 14418 312044 14424
rect 310796 9104 310848 9110
rect 310796 9046 310848 9052
rect 310704 9036 310756 9042
rect 310704 8978 310756 8984
rect 312096 7886 312124 316006
rect 312084 7880 312136 7886
rect 312084 7822 312136 7828
rect 310612 7812 310664 7818
rect 310612 7754 310664 7760
rect 313292 6186 313320 330482
rect 313384 7954 313412 338014
rect 313752 316034 313780 338014
rect 314120 330546 314148 338014
rect 314108 330540 314160 330546
rect 314108 330482 314160 330488
rect 314752 327208 314804 327214
rect 314752 327150 314804 327156
rect 313476 316006 313780 316034
rect 313476 10334 313504 316006
rect 313464 10328 313516 10334
rect 313464 10270 313516 10276
rect 314764 8090 314792 327150
rect 314752 8084 314804 8090
rect 314752 8026 314804 8032
rect 314856 8022 314884 338014
rect 314948 338014 315100 338042
rect 315224 338014 315468 338042
rect 315592 338014 315836 338042
rect 316052 338014 316204 338042
rect 316328 338014 316572 338042
rect 316696 338014 316940 338042
rect 317064 338014 317308 338042
rect 317524 338014 317676 338042
rect 317800 338014 318044 338042
rect 318168 338014 318412 338042
rect 318536 338014 318780 338042
rect 318996 338014 319148 338042
rect 319272 338014 319424 338042
rect 319548 338014 319792 338042
rect 319916 338014 320160 338042
rect 320284 338014 320528 338042
rect 320652 338014 320896 338042
rect 321020 338014 321264 338042
rect 321572 338014 321632 338042
rect 321756 338014 322000 338042
rect 322124 338014 322368 338042
rect 322492 338014 322736 338042
rect 323044 338014 323104 338042
rect 323228 338014 323472 338042
rect 323596 338014 323840 338042
rect 323964 338014 324208 338042
rect 324516 338014 324576 338042
rect 324700 338014 324944 338042
rect 325068 338014 325312 338042
rect 325436 338014 325680 338042
rect 325988 338014 326048 338042
rect 326172 338014 326416 338042
rect 326540 338014 326784 338042
rect 327092 338014 327152 338042
rect 327276 338014 327520 338042
rect 327644 338014 327888 338042
rect 328012 338014 328256 338042
rect 328472 338014 328624 338042
rect 328748 338014 328992 338042
rect 329116 338014 329360 338042
rect 329484 338014 329728 338042
rect 330036 338014 330096 338042
rect 330220 338014 330464 338042
rect 330588 338014 330832 338042
rect 330956 338014 331108 338042
rect 331476 338014 331628 338042
rect 314948 335646 314976 338014
rect 315224 335986 315252 338014
rect 315212 335980 315264 335986
rect 315212 335922 315264 335928
rect 314936 335640 314988 335646
rect 314936 335582 314988 335588
rect 315592 327214 315620 338014
rect 316052 336054 316080 338014
rect 316328 336682 316356 338014
rect 316144 336654 316356 336682
rect 316040 336048 316092 336054
rect 316040 335990 316092 335996
rect 315580 327208 315632 327214
rect 315580 327150 315632 327156
rect 316144 10402 316172 336654
rect 316696 336546 316724 338014
rect 316236 336518 316724 336546
rect 316132 10396 316184 10402
rect 316132 10338 316184 10344
rect 316236 8158 316264 336518
rect 317064 336190 317092 338014
rect 317052 336184 317104 336190
rect 317052 336126 317104 336132
rect 316684 336048 316736 336054
rect 316684 335990 316736 335996
rect 316224 8152 316276 8158
rect 316224 8094 316276 8100
rect 314844 8016 314896 8022
rect 314844 7958 314896 7964
rect 313372 7948 313424 7954
rect 313372 7890 313424 7896
rect 316696 6390 316724 335990
rect 317524 10470 317552 338014
rect 317604 330540 317656 330546
rect 317604 330482 317656 330488
rect 317616 10538 317644 330482
rect 317800 316034 317828 338014
rect 318168 336122 318196 338014
rect 318156 336116 318208 336122
rect 318156 336058 318208 336064
rect 318536 330546 318564 338014
rect 318524 330540 318576 330546
rect 318524 330482 318576 330488
rect 318892 330540 318944 330546
rect 318892 330482 318944 330488
rect 317708 316006 317828 316034
rect 317604 10532 317656 10538
rect 317604 10474 317656 10480
rect 317512 10464 317564 10470
rect 317512 10406 317564 10412
rect 316684 6384 316736 6390
rect 316684 6326 316736 6332
rect 317708 6254 317736 316006
rect 317696 6248 317748 6254
rect 317696 6190 317748 6196
rect 313280 6180 313332 6186
rect 313280 6122 313332 6128
rect 318904 5098 318932 330482
rect 318892 5092 318944 5098
rect 318892 5034 318944 5040
rect 310520 5024 310572 5030
rect 310520 4966 310572 4972
rect 309140 4956 309192 4962
rect 309140 4898 309192 4904
rect 307760 4888 307812 4894
rect 307760 4830 307812 4836
rect 306472 4548 306524 4554
rect 306472 4490 306524 4496
rect 309048 4140 309100 4146
rect 309048 4082 309100 4088
rect 307944 4072 307996 4078
rect 307944 4014 307996 4020
rect 305552 4004 305604 4010
rect 305552 3946 305604 3952
rect 304356 3392 304408 3398
rect 304356 3334 304408 3340
rect 304908 3392 304960 3398
rect 304908 3334 304960 3340
rect 304368 480 304396 3334
rect 305564 480 305592 3946
rect 306748 3392 306800 3398
rect 306748 3334 306800 3340
rect 306760 480 306788 3334
rect 307956 480 307984 4014
rect 309060 480 309088 4082
rect 318996 3466 319024 338014
rect 319272 336258 319300 338014
rect 319260 336252 319312 336258
rect 319260 336194 319312 336200
rect 319548 330546 319576 338014
rect 319916 336394 319944 338014
rect 319904 336388 319956 336394
rect 319904 336330 319956 336336
rect 319536 330540 319588 330546
rect 319536 330482 319588 330488
rect 320180 330540 320232 330546
rect 320180 330482 320232 330488
rect 320192 3534 320220 330482
rect 320180 3528 320232 3534
rect 320180 3470 320232 3476
rect 318984 3460 319036 3466
rect 318984 3402 319036 3408
rect 319720 3460 319772 3466
rect 319720 3402 319772 3408
rect 310244 3324 310296 3330
rect 310244 3266 310296 3272
rect 310256 480 310284 3266
rect 311440 3256 311492 3262
rect 311440 3198 311492 3204
rect 311452 480 311480 3198
rect 312636 3188 312688 3194
rect 312636 3130 312688 3136
rect 312648 480 312676 3130
rect 313832 3120 313884 3126
rect 313832 3062 313884 3068
rect 313844 480 313872 3062
rect 315028 3052 315080 3058
rect 315028 2994 315080 3000
rect 315040 480 315068 2994
rect 317328 2984 317380 2990
rect 317328 2926 317380 2932
rect 316224 2848 316276 2854
rect 316224 2790 316276 2796
rect 316236 480 316264 2790
rect 317340 480 317368 2926
rect 318524 2916 318576 2922
rect 318524 2858 318576 2864
rect 318536 480 318564 2858
rect 319732 480 319760 3402
rect 320284 3369 320312 338014
rect 320652 316034 320680 338014
rect 321020 330546 321048 338014
rect 321572 336326 321600 338014
rect 321560 336320 321612 336326
rect 321560 336262 321612 336268
rect 321008 330540 321060 330546
rect 321008 330482 321060 330488
rect 321652 330540 321704 330546
rect 321652 330482 321704 330488
rect 320376 316006 320680 316034
rect 320376 5166 320404 316006
rect 320364 5160 320416 5166
rect 320364 5102 320416 5108
rect 320916 3868 320968 3874
rect 320916 3810 320968 3816
rect 320270 3360 320326 3369
rect 320270 3295 320326 3304
rect 320928 480 320956 3810
rect 321664 3505 321692 330482
rect 321756 4486 321784 338014
rect 322124 330546 322152 338014
rect 322112 330540 322164 330546
rect 322112 330482 322164 330488
rect 322492 316034 322520 338014
rect 321848 316006 322520 316034
rect 321744 4480 321796 4486
rect 321744 4422 321796 4428
rect 321848 3602 321876 316006
rect 323044 4418 323072 338014
rect 323124 330540 323176 330546
rect 323124 330482 323176 330488
rect 323032 4412 323084 4418
rect 323032 4354 323084 4360
rect 323136 4350 323164 330482
rect 323124 4344 323176 4350
rect 323124 4286 323176 4292
rect 323228 3670 323256 338014
rect 323596 336462 323624 338014
rect 323584 336456 323636 336462
rect 323584 336398 323636 336404
rect 323964 330546 323992 338014
rect 323952 330540 324004 330546
rect 323952 330482 324004 330488
rect 324320 330540 324372 330546
rect 324320 330482 324372 330488
rect 324332 4026 324360 330482
rect 324412 330472 324464 330478
rect 324412 330414 324464 330420
rect 324240 3998 324360 4026
rect 324240 3670 324268 3998
rect 324424 3924 324452 330414
rect 324332 3896 324452 3924
rect 324332 3806 324360 3896
rect 324320 3800 324372 3806
rect 324320 3742 324372 3748
rect 324412 3800 324464 3806
rect 324412 3742 324464 3748
rect 323216 3664 323268 3670
rect 323216 3606 323268 3612
rect 324228 3664 324280 3670
rect 324228 3606 324280 3612
rect 321836 3596 321888 3602
rect 321836 3538 321888 3544
rect 323400 3596 323452 3602
rect 323400 3538 323452 3544
rect 322112 3528 322164 3534
rect 321650 3496 321706 3505
rect 322112 3470 322164 3476
rect 321650 3431 321706 3440
rect 322124 480 322152 3470
rect 323412 1850 323440 3538
rect 323320 1822 323440 1850
rect 323320 480 323348 1822
rect 324424 480 324452 3742
rect 324516 3641 324544 338014
rect 324700 330546 324728 338014
rect 324688 330540 324740 330546
rect 324688 330482 324740 330488
rect 325068 316034 325096 338014
rect 325436 330478 325464 338014
rect 325792 330540 325844 330546
rect 325792 330482 325844 330488
rect 325424 330472 325476 330478
rect 325424 330414 325476 330420
rect 324608 316006 325096 316034
rect 324608 4282 324636 316006
rect 324596 4276 324648 4282
rect 324596 4218 324648 4224
rect 325804 3942 325832 330482
rect 325792 3936 325844 3942
rect 325792 3878 325844 3884
rect 325988 3777 326016 338014
rect 326172 336598 326200 338014
rect 326160 336592 326212 336598
rect 326160 336534 326212 336540
rect 326540 330546 326568 338014
rect 327092 336530 327120 338014
rect 327080 336524 327132 336530
rect 327080 336466 327132 336472
rect 327276 336054 327304 338014
rect 327644 336818 327672 338014
rect 327552 336790 327672 336818
rect 327552 336666 327580 336790
rect 328012 336682 328040 338014
rect 327540 336660 327592 336666
rect 327540 336602 327592 336608
rect 327644 336654 328040 336682
rect 327264 336048 327316 336054
rect 327264 335990 327316 335996
rect 326528 330540 326580 330546
rect 326528 330482 326580 330488
rect 327644 316034 327672 336654
rect 328472 336258 328500 338014
rect 328748 336954 328776 338014
rect 328564 336926 328776 336954
rect 328564 336734 328592 336926
rect 329116 336818 329144 338014
rect 328656 336790 329144 336818
rect 328552 336728 328604 336734
rect 328552 336670 328604 336676
rect 327724 336252 327776 336258
rect 327724 336194 327776 336200
rect 328460 336252 328512 336258
rect 328460 336194 328512 336200
rect 327276 316006 327672 316034
rect 327276 3806 327304 316006
rect 327736 6322 327764 336194
rect 328368 336048 328420 336054
rect 328368 335990 328420 335996
rect 327724 6316 327776 6322
rect 327724 6258 327776 6264
rect 327264 3800 327316 3806
rect 325974 3768 326030 3777
rect 327264 3742 327316 3748
rect 325974 3703 326030 3712
rect 326804 3732 326856 3738
rect 326804 3674 326856 3680
rect 325608 3664 325660 3670
rect 324502 3632 324558 3641
rect 325608 3606 325660 3612
rect 324502 3567 324558 3576
rect 325620 480 325648 3606
rect 326816 480 326844 3674
rect 328012 598 328224 626
rect 328012 480 328040 598
rect 328196 490 328224 598
rect 328380 490 328408 335990
rect 328656 316034 328684 336790
rect 329484 336682 329512 338014
rect 329024 336654 329512 336682
rect 329024 316034 329052 336654
rect 329104 336524 329156 336530
rect 329104 336466 329156 336472
rect 328564 316006 328684 316034
rect 328748 316006 329052 316034
rect 328564 4010 328592 316006
rect 328552 4004 328604 4010
rect 328552 3946 328604 3952
rect 328748 3398 328776 316006
rect 329116 3874 329144 336466
rect 329932 330540 329984 330546
rect 329932 330482 329984 330488
rect 329840 328092 329892 328098
rect 329840 328034 329892 328040
rect 329196 4004 329248 4010
rect 329196 3946 329248 3952
rect 329104 3868 329156 3874
rect 329104 3810 329156 3816
rect 328736 3392 328788 3398
rect 328736 3334 328788 3340
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 328196 462 328408 490
rect 329208 480 329236 3946
rect 329852 3330 329880 328034
rect 329840 3324 329892 3330
rect 329840 3266 329892 3272
rect 329944 3262 329972 330482
rect 330036 4078 330064 338014
rect 330220 316034 330248 338014
rect 330588 328098 330616 338014
rect 330956 330546 330984 338014
rect 331600 330818 331628 338014
rect 331692 338014 331844 338042
rect 331968 338014 332212 338042
rect 332336 338014 332580 338042
rect 332704 338014 332948 338042
rect 333072 338014 333316 338042
rect 333440 338014 333684 338042
rect 333992 338014 334052 338042
rect 334176 338014 334420 338042
rect 334544 338014 334788 338042
rect 334912 338014 335156 338042
rect 331588 330812 331640 330818
rect 331588 330754 331640 330760
rect 331692 330698 331720 338014
rect 331416 330670 331720 330698
rect 330944 330540 330996 330546
rect 330944 330482 330996 330488
rect 331312 330472 331364 330478
rect 331312 330414 331364 330420
rect 330576 328092 330628 328098
rect 330576 328034 330628 328040
rect 330128 316006 330248 316034
rect 330128 4146 330156 316006
rect 330116 4140 330168 4146
rect 330116 4082 330168 4088
rect 330024 4072 330076 4078
rect 330024 4014 330076 4020
rect 331220 3800 331272 3806
rect 331220 3742 331272 3748
rect 329932 3256 329984 3262
rect 329932 3198 329984 3204
rect 330392 3188 330444 3194
rect 330392 3130 330444 3136
rect 330404 480 330432 3130
rect 331232 3058 331260 3742
rect 331220 3052 331272 3058
rect 331220 2994 331272 3000
rect 331324 2854 331352 330414
rect 331416 3126 331444 330670
rect 331588 330608 331640 330614
rect 331588 330550 331640 330556
rect 331496 330540 331548 330546
rect 331496 330482 331548 330488
rect 331508 3806 331536 330482
rect 331496 3800 331548 3806
rect 331496 3742 331548 3748
rect 331600 3618 331628 330550
rect 331968 330546 331996 338014
rect 331956 330540 332008 330546
rect 331956 330482 332008 330488
rect 332336 330478 332364 338014
rect 332508 335368 332560 335374
rect 332508 335310 332560 335316
rect 332324 330472 332376 330478
rect 332324 330414 332376 330420
rect 331508 3590 331628 3618
rect 331508 3262 331536 3590
rect 332520 3534 332548 335310
rect 332600 330540 332652 330546
rect 332600 330482 332652 330488
rect 331588 3528 331640 3534
rect 331588 3470 331640 3476
rect 332508 3528 332560 3534
rect 332508 3470 332560 3476
rect 331496 3256 331548 3262
rect 331496 3198 331548 3204
rect 331404 3120 331456 3126
rect 331404 3062 331456 3068
rect 331312 2848 331364 2854
rect 331312 2790 331364 2796
rect 331600 480 331628 3470
rect 332612 3466 332640 330482
rect 332704 6914 332732 338014
rect 333072 316034 333100 338014
rect 333244 335912 333296 335918
rect 333244 335854 333296 335860
rect 332796 316006 333100 316034
rect 332796 16574 332824 316006
rect 332796 16546 332916 16574
rect 332704 6886 332824 6914
rect 332692 4140 332744 4146
rect 332692 4082 332744 4088
rect 332600 3460 332652 3466
rect 332600 3402 332652 3408
rect 332704 480 332732 4082
rect 332796 2990 332824 6886
rect 332784 2984 332836 2990
rect 332784 2926 332836 2932
rect 332888 2922 332916 16546
rect 333256 3194 333284 335854
rect 333440 330546 333468 338014
rect 333992 336530 334020 338014
rect 333980 336524 334032 336530
rect 333980 336466 334032 336472
rect 333428 330540 333480 330546
rect 333428 330482 333480 330488
rect 334072 330540 334124 330546
rect 334072 330482 334124 330488
rect 333888 3868 333940 3874
rect 333888 3810 333940 3816
rect 333244 3188 333296 3194
rect 333244 3130 333296 3136
rect 332876 2916 332928 2922
rect 332876 2858 332928 2864
rect 333900 480 333928 3810
rect 334084 3602 334112 330482
rect 334072 3596 334124 3602
rect 334072 3538 334124 3544
rect 334176 3398 334204 338014
rect 334544 330546 334572 338014
rect 334532 330540 334584 330546
rect 334532 330482 334584 330488
rect 334912 316034 334940 338014
rect 335510 337770 335538 338028
rect 335648 338014 335892 338042
rect 336016 338014 336260 338042
rect 336384 338014 336628 338042
rect 336752 338014 336996 338042
rect 337120 338014 337364 338042
rect 337488 338014 337732 338042
rect 337856 338014 338100 338042
rect 338316 338014 338468 338042
rect 338592 338014 338836 338042
rect 338960 338014 339204 338042
rect 335510 337742 335584 337770
rect 335452 330540 335504 330546
rect 335452 330482 335504 330488
rect 334268 316006 334940 316034
rect 334268 3942 334296 316006
rect 335464 4010 335492 330482
rect 335452 4004 335504 4010
rect 335452 3946 335504 3952
rect 334256 3936 334308 3942
rect 334256 3878 334308 3884
rect 335556 3670 335584 337742
rect 335648 3738 335676 338014
rect 336016 336054 336044 338014
rect 336004 336048 336056 336054
rect 336004 335990 336056 335996
rect 336004 335844 336056 335850
rect 336004 335786 336056 335792
rect 336016 4146 336044 335786
rect 336384 330546 336412 338014
rect 336752 335918 336780 338014
rect 336740 335912 336792 335918
rect 336740 335854 336792 335860
rect 337120 335374 337148 338014
rect 337488 335850 337516 338014
rect 337476 335844 337528 335850
rect 337476 335786 337528 335792
rect 337108 335368 337160 335374
rect 337108 335310 337160 335316
rect 336372 330540 336424 330546
rect 336372 330482 336424 330488
rect 337856 316034 337884 338014
rect 338120 330540 338172 330546
rect 338120 330482 338172 330488
rect 336936 316006 337884 316034
rect 336004 4140 336056 4146
rect 336004 4082 336056 4088
rect 336936 3874 336964 316006
rect 336924 3868 336976 3874
rect 336924 3810 336976 3816
rect 335636 3732 335688 3738
rect 335636 3674 335688 3680
rect 335544 3664 335596 3670
rect 335544 3606 335596 3612
rect 338132 3534 338160 330482
rect 338212 330472 338264 330478
rect 338212 330414 338264 330420
rect 336280 3528 336332 3534
rect 336280 3470 336332 3476
rect 338120 3528 338172 3534
rect 338120 3470 338172 3476
rect 335084 3460 335136 3466
rect 335084 3402 335136 3408
rect 334164 3392 334216 3398
rect 334164 3334 334216 3340
rect 335096 480 335124 3402
rect 336292 480 336320 3470
rect 338224 3058 338252 330414
rect 338316 3466 338344 338014
rect 338592 330546 338620 338014
rect 338580 330540 338632 330546
rect 338580 330482 338632 330488
rect 338960 330478 338988 338014
rect 339558 337770 339586 338028
rect 339788 338014 339940 338042
rect 340308 338014 340552 338042
rect 340676 338014 340828 338042
rect 341044 338014 341288 338042
rect 341412 338014 341656 338042
rect 341780 338014 342024 338042
rect 339558 337742 339632 337770
rect 339500 336728 339552 336734
rect 339500 336670 339552 336676
rect 338948 330472 339000 330478
rect 338948 330414 339000 330420
rect 338304 3460 338356 3466
rect 338304 3402 338356 3408
rect 338672 3120 338724 3126
rect 338672 3062 338724 3068
rect 337476 3052 337528 3058
rect 337476 2994 337528 3000
rect 338212 3052 338264 3058
rect 338212 2994 338264 3000
rect 337488 480 337516 2994
rect 338684 480 338712 3062
rect 339512 490 339540 336670
rect 339604 3126 339632 337742
rect 339788 336734 339816 338014
rect 339776 336728 339828 336734
rect 339776 336670 339828 336676
rect 340524 335354 340552 338014
rect 340800 336682 340828 338014
rect 340800 336654 341196 336682
rect 341260 336666 341288 338014
rect 340524 335326 340828 335354
rect 340800 3482 340828 335326
rect 341168 16574 341196 336654
rect 341248 336660 341300 336666
rect 341248 336602 341300 336608
rect 341628 336258 341656 338014
rect 341616 336252 341668 336258
rect 341616 336194 341668 336200
rect 341996 335442 342024 338014
rect 342088 338014 342148 338042
rect 342516 338014 342760 338042
rect 342884 338014 343036 338042
rect 343160 338014 343404 338042
rect 341984 335436 342036 335442
rect 341984 335378 342036 335384
rect 341168 16546 342024 16574
rect 340800 3454 341012 3482
rect 339592 3120 339644 3126
rect 339592 3062 339644 3068
rect 339696 598 339908 626
rect 339696 490 339724 598
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339512 462 339724 490
rect 339880 480 339908 598
rect 340984 480 341012 3454
rect 341996 3074 342024 16546
rect 342088 3602 342116 338014
rect 342732 336734 342760 338014
rect 342720 336728 342772 336734
rect 342720 336670 342772 336676
rect 342444 336660 342496 336666
rect 342444 336602 342496 336608
rect 342168 336252 342220 336258
rect 342168 336194 342220 336200
rect 342076 3596 342128 3602
rect 342076 3538 342128 3544
rect 342180 3194 342208 336194
rect 342456 16574 342484 336602
rect 343008 325694 343036 338014
rect 343376 330426 343404 338014
rect 343514 337770 343542 338028
rect 343896 338014 344140 338042
rect 344264 338014 344508 338042
rect 344632 338014 344876 338042
rect 343514 337742 343588 337770
rect 343560 336734 343588 337742
rect 343456 336728 343508 336734
rect 343456 336670 343508 336676
rect 343548 336728 343600 336734
rect 343548 336670 343600 336676
rect 343468 330562 343496 336670
rect 344112 336122 344140 338014
rect 344284 336728 344336 336734
rect 344284 336670 344336 336676
rect 344100 336116 344152 336122
rect 344100 336058 344152 336064
rect 343468 330534 343588 330562
rect 343376 330398 343496 330426
rect 343008 325666 343404 325694
rect 342456 16546 342944 16574
rect 342168 3188 342220 3194
rect 342168 3130 342220 3136
rect 341996 3046 342208 3074
rect 342180 480 342208 3046
rect 342916 490 342944 16546
rect 343376 4010 343404 325666
rect 343468 4146 343496 330398
rect 343456 4140 343508 4146
rect 343456 4082 343508 4088
rect 343560 4078 343588 330534
rect 343548 4072 343600 4078
rect 343548 4014 343600 4020
rect 343364 4004 343416 4010
rect 343364 3946 343416 3952
rect 344296 3942 344324 336670
rect 344480 335578 344508 338014
rect 344848 336054 344876 338014
rect 344940 338014 345000 338042
rect 345368 338014 345612 338042
rect 345736 338014 345980 338042
rect 346104 338014 346348 338042
rect 346472 338014 346716 338042
rect 346840 338014 347084 338042
rect 347208 338014 347452 338042
rect 347576 338014 347728 338042
rect 347944 338014 348188 338042
rect 348312 338014 348556 338042
rect 348680 338014 348924 338042
rect 344836 336048 344888 336054
rect 344836 335990 344888 335996
rect 344468 335572 344520 335578
rect 344468 335514 344520 335520
rect 344940 335374 344968 338014
rect 345584 336598 345612 338014
rect 345572 336592 345624 336598
rect 345572 336534 345624 336540
rect 345664 336116 345716 336122
rect 345664 336058 345716 336064
rect 345204 335436 345256 335442
rect 345204 335378 345256 335384
rect 344928 335368 344980 335374
rect 344928 335310 344980 335316
rect 345216 16574 345244 335378
rect 345216 16546 345336 16574
rect 344284 3936 344336 3942
rect 344284 3878 344336 3884
rect 344560 3188 344612 3194
rect 344560 3130 344612 3136
rect 343192 598 343404 626
rect 343192 490 343220 598
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 462 343220 490
rect 343376 480 343404 598
rect 344572 480 344600 3130
rect 345308 490 345336 16546
rect 345676 3534 345704 336058
rect 345756 335368 345808 335374
rect 345756 335310 345808 335316
rect 345768 3874 345796 335310
rect 345952 325694 345980 338014
rect 346320 335986 346348 338014
rect 346688 336258 346716 338014
rect 347056 336734 347084 338014
rect 347044 336728 347096 336734
rect 347044 336670 347096 336676
rect 347424 336462 347452 338014
rect 347596 336728 347648 336734
rect 347596 336670 347648 336676
rect 347412 336456 347464 336462
rect 347412 336398 347464 336404
rect 346676 336252 346728 336258
rect 346676 336194 346728 336200
rect 346308 335980 346360 335986
rect 346308 335922 346360 335928
rect 347136 335980 347188 335986
rect 347136 335922 347188 335928
rect 346952 335572 347004 335578
rect 346952 335514 347004 335520
rect 346964 325694 346992 335514
rect 345952 325666 346348 325694
rect 346964 325666 347084 325694
rect 345756 3868 345808 3874
rect 345756 3810 345808 3816
rect 346320 3806 346348 325666
rect 346308 3800 346360 3806
rect 346308 3742 346360 3748
rect 346952 3596 347004 3602
rect 346952 3538 347004 3544
rect 345664 3528 345716 3534
rect 345664 3470 345716 3476
rect 345584 598 345796 626
rect 345584 490 345612 598
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345308 462 345612 490
rect 345768 480 345796 598
rect 346964 480 346992 3538
rect 347056 3194 347084 325666
rect 347148 3670 347176 335922
rect 347608 3738 347636 336670
rect 347700 336394 347728 338014
rect 347688 336388 347740 336394
rect 347688 336330 347740 336336
rect 347688 336252 347740 336258
rect 347688 336194 347740 336200
rect 347596 3732 347648 3738
rect 347596 3674 347648 3680
rect 347136 3664 347188 3670
rect 347136 3606 347188 3612
rect 347700 3602 347728 336194
rect 348160 336122 348188 338014
rect 348528 336530 348556 338014
rect 348516 336524 348568 336530
rect 348516 336466 348568 336472
rect 348424 336388 348476 336394
rect 348424 336330 348476 336336
rect 348148 336116 348200 336122
rect 348148 336058 348200 336064
rect 348056 4072 348108 4078
rect 348056 4014 348108 4020
rect 347688 3596 347740 3602
rect 347688 3538 347740 3544
rect 347044 3188 347096 3194
rect 347044 3130 347096 3136
rect 348068 480 348096 4014
rect 348436 3058 348464 336330
rect 348896 336326 348924 338014
rect 348988 338014 349048 338042
rect 349416 338014 349660 338042
rect 349784 338014 350028 338042
rect 348884 336320 348936 336326
rect 348884 336262 348936 336268
rect 348516 336048 348568 336054
rect 348516 335990 348568 335996
rect 348528 3398 348556 335990
rect 348988 3466 349016 338014
rect 349632 336666 349660 338014
rect 349620 336660 349672 336666
rect 349620 336602 349672 336608
rect 349804 336592 349856 336598
rect 349804 336534 349856 336540
rect 349068 336116 349120 336122
rect 349068 336058 349120 336064
rect 348976 3460 349028 3466
rect 348976 3402 349028 3408
rect 348516 3392 348568 3398
rect 348516 3334 348568 3340
rect 349080 3262 349108 336058
rect 349252 4004 349304 4010
rect 349252 3946 349304 3952
rect 349068 3256 349120 3262
rect 349068 3198 349120 3204
rect 348424 3052 348476 3058
rect 348424 2994 348476 3000
rect 349264 480 349292 3946
rect 349816 3126 349844 336534
rect 350000 330546 350028 338014
rect 350092 338014 350152 338042
rect 350276 338014 350520 338042
rect 350888 338014 351132 338042
rect 351256 338014 351500 338042
rect 351624 338014 351776 338042
rect 351992 338014 352236 338042
rect 352360 338014 352604 338042
rect 352728 338014 352972 338042
rect 350092 335442 350120 338014
rect 350080 335436 350132 335442
rect 350080 335378 350132 335384
rect 349988 330540 350040 330546
rect 349988 330482 350040 330488
rect 350276 4486 350304 338014
rect 351104 336122 351132 338014
rect 351472 336190 351500 338014
rect 351460 336184 351512 336190
rect 351460 336126 351512 336132
rect 351092 336116 351144 336122
rect 351092 336058 351144 336064
rect 350356 335436 350408 335442
rect 350356 335378 350408 335384
rect 350264 4480 350316 4486
rect 350264 4422 350316 4428
rect 350368 4078 350396 335378
rect 350448 330540 350500 330546
rect 350448 330482 350500 330488
rect 350460 4298 350488 330482
rect 351748 4554 351776 338014
rect 352208 336258 352236 338014
rect 352196 336252 352248 336258
rect 352196 336194 352248 336200
rect 352576 336122 352604 338014
rect 351828 336116 351880 336122
rect 351828 336058 351880 336064
rect 352564 336116 352616 336122
rect 352564 336058 352616 336064
rect 351736 4548 351788 4554
rect 351736 4490 351788 4496
rect 350460 4270 350580 4298
rect 350448 4140 350500 4146
rect 350448 4082 350500 4088
rect 350356 4072 350408 4078
rect 350356 4014 350408 4020
rect 349804 3120 349856 3126
rect 349804 3062 349856 3068
rect 350460 480 350488 4082
rect 350552 3330 350580 4270
rect 351840 4146 351868 336058
rect 352944 335578 352972 338014
rect 353036 338014 353096 338042
rect 353464 338014 353708 338042
rect 353832 338014 354076 338042
rect 354200 338014 354444 338042
rect 352932 335572 352984 335578
rect 352932 335514 352984 335520
rect 353036 8974 353064 338014
rect 353208 336116 353260 336122
rect 353208 336058 353260 336064
rect 353116 335572 353168 335578
rect 353116 335514 353168 335520
rect 353024 8968 353076 8974
rect 353024 8910 353076 8916
rect 353128 4622 353156 335514
rect 353116 4616 353168 4622
rect 353116 4558 353168 4564
rect 351828 4140 351880 4146
rect 351828 4082 351880 4088
rect 353220 4010 353248 336058
rect 353680 336054 353708 338014
rect 354048 336734 354076 338014
rect 354036 336728 354088 336734
rect 354036 336670 354088 336676
rect 353944 336660 353996 336666
rect 353944 336602 353996 336608
rect 353668 336048 353720 336054
rect 353668 335990 353720 335996
rect 353956 9042 353984 336602
rect 354416 336394 354444 338014
rect 354554 337770 354582 338028
rect 354936 338014 355088 338042
rect 355212 338014 355456 338042
rect 355580 338014 355732 338042
rect 354554 337742 354628 337770
rect 354496 336728 354548 336734
rect 354496 336670 354548 336676
rect 354404 336388 354456 336394
rect 354404 336330 354456 336336
rect 353944 9036 353996 9042
rect 353944 8978 353996 8984
rect 354508 4690 354536 336670
rect 354496 4684 354548 4690
rect 354496 4626 354548 4632
rect 353208 4004 353260 4010
rect 353208 3946 353260 3952
rect 354600 3942 354628 337742
rect 355060 336734 355088 338014
rect 355048 336728 355100 336734
rect 355048 336670 355100 336676
rect 355428 335374 355456 338014
rect 355704 336666 355732 338014
rect 355888 338014 355948 338042
rect 356316 338014 356560 338042
rect 356684 338014 356928 338042
rect 357052 338014 357296 338042
rect 355784 336728 355836 336734
rect 355784 336670 355836 336676
rect 355692 336660 355744 336666
rect 355692 336602 355744 336608
rect 355416 335368 355468 335374
rect 355416 335310 355468 335316
rect 355796 4758 355824 336670
rect 355888 5506 355916 338014
rect 356532 336734 356560 338014
rect 356520 336728 356572 336734
rect 356520 336670 356572 336676
rect 355968 336660 356020 336666
rect 355968 336602 356020 336608
rect 355876 5500 355928 5506
rect 355876 5442 355928 5448
rect 355784 4752 355836 4758
rect 355784 4694 355836 4700
rect 351644 3936 351696 3942
rect 351644 3878 351696 3884
rect 354588 3936 354640 3942
rect 354588 3878 354640 3884
rect 350540 3324 350592 3330
rect 350540 3266 350592 3272
rect 351656 480 351684 3878
rect 352840 3528 352892 3534
rect 352840 3470 352892 3476
rect 352852 480 352880 3470
rect 355232 3392 355284 3398
rect 355232 3334 355284 3340
rect 354036 3188 354088 3194
rect 354036 3130 354088 3136
rect 354048 480 354076 3130
rect 355244 480 355272 3334
rect 355980 2990 356008 336602
rect 356900 335986 356928 338014
rect 357164 336728 357216 336734
rect 357164 336670 357216 336676
rect 356888 335980 356940 335986
rect 356888 335922 356940 335928
rect 357176 10334 357204 336670
rect 357164 10328 357216 10334
rect 357164 10270 357216 10276
rect 357268 5438 357296 338014
rect 357360 338014 357420 338042
rect 357788 338014 358032 338042
rect 358156 338014 358400 338042
rect 358524 338014 358676 338042
rect 358892 338014 359136 338042
rect 359260 338014 359504 338042
rect 359628 338014 359872 338042
rect 359996 338014 360148 338042
rect 360364 338014 360608 338042
rect 360732 338014 360976 338042
rect 357360 336138 357388 338014
rect 358004 336734 358032 338014
rect 357992 336728 358044 336734
rect 357992 336670 358044 336676
rect 358084 336184 358136 336190
rect 357360 336110 357480 336138
rect 358084 336126 358136 336132
rect 357348 335980 357400 335986
rect 357348 335922 357400 335928
rect 357256 5432 357308 5438
rect 357256 5374 357308 5380
rect 357360 3874 357388 335922
rect 357452 335442 357480 336110
rect 357440 335436 357492 335442
rect 357440 335378 357492 335384
rect 356336 3868 356388 3874
rect 356336 3810 356388 3816
rect 357348 3868 357400 3874
rect 357348 3810 357400 3816
rect 355968 2984 356020 2990
rect 355968 2926 356020 2932
rect 356348 480 356376 3810
rect 358096 3738 358124 336126
rect 358372 335354 358400 338014
rect 358372 335326 358584 335354
rect 358556 5302 358584 335326
rect 358648 5370 358676 338014
rect 358728 336728 358780 336734
rect 358728 336670 358780 336676
rect 358636 5364 358688 5370
rect 358636 5306 358688 5312
rect 358544 5296 358596 5302
rect 358544 5238 358596 5244
rect 358740 3806 358768 336670
rect 359108 336666 359136 338014
rect 359476 336734 359504 338014
rect 359464 336728 359516 336734
rect 359464 336670 359516 336676
rect 359096 336660 359148 336666
rect 359096 336602 359148 336608
rect 359844 5166 359872 338014
rect 359924 336728 359976 336734
rect 359924 336670 359976 336676
rect 359936 5234 359964 336670
rect 360016 336660 360068 336666
rect 360016 336602 360068 336608
rect 359924 5228 359976 5234
rect 359924 5170 359976 5176
rect 359832 5160 359884 5166
rect 359832 5102 359884 5108
rect 358728 3800 358780 3806
rect 358728 3742 358780 3748
rect 358084 3732 358136 3738
rect 358084 3674 358136 3680
rect 360028 3670 360056 336602
rect 358728 3664 358780 3670
rect 358728 3606 358780 3612
rect 360016 3664 360068 3670
rect 360016 3606 360068 3612
rect 357532 3120 357584 3126
rect 357532 3062 357584 3068
rect 357544 480 357572 3062
rect 358740 480 358768 3606
rect 360120 3602 360148 338014
rect 360580 335714 360608 338014
rect 360948 336734 360976 338014
rect 361040 338014 361100 338042
rect 361224 338014 361468 338042
rect 361836 338014 362080 338042
rect 362204 338014 362448 338042
rect 362572 338014 362816 338042
rect 360936 336728 360988 336734
rect 360936 336670 360988 336676
rect 361040 335850 361068 338014
rect 361028 335844 361080 335850
rect 361028 335786 361080 335792
rect 360568 335708 360620 335714
rect 360568 335650 360620 335656
rect 361224 4894 361252 338014
rect 361396 336728 361448 336734
rect 361396 336670 361448 336676
rect 361304 335708 361356 335714
rect 361304 335650 361356 335656
rect 361316 5098 361344 335650
rect 361304 5092 361356 5098
rect 361304 5034 361356 5040
rect 361408 5030 361436 336670
rect 362052 336666 362080 338014
rect 362040 336660 362092 336666
rect 362040 336602 362092 336608
rect 361488 335844 361540 335850
rect 361488 335786 361540 335792
rect 361396 5024 361448 5030
rect 361396 4966 361448 4972
rect 361212 4888 361264 4894
rect 361212 4830 361264 4836
rect 359924 3596 359976 3602
rect 359924 3538 359976 3544
rect 360108 3596 360160 3602
rect 360108 3538 360160 3544
rect 359936 480 359964 3538
rect 361500 3534 361528 335786
rect 362420 330546 362448 338014
rect 362592 336728 362644 336734
rect 362592 336670 362644 336676
rect 362408 330540 362460 330546
rect 362408 330482 362460 330488
rect 362604 7070 362632 336670
rect 362684 336660 362736 336666
rect 362684 336602 362736 336608
rect 362592 7064 362644 7070
rect 362592 7006 362644 7012
rect 362696 4962 362724 336602
rect 362684 4956 362736 4962
rect 362684 4898 362736 4904
rect 362788 4826 362816 338014
rect 362880 338014 362940 338042
rect 363308 338014 363552 338042
rect 363676 338014 363920 338042
rect 364044 338014 364196 338042
rect 364412 338014 364656 338042
rect 364780 338014 365024 338042
rect 365148 338014 365392 338042
rect 365516 338014 365668 338042
rect 365884 338014 366128 338042
rect 366252 338014 366496 338042
rect 366620 338014 366864 338042
rect 362880 336734 362908 338014
rect 363524 336734 363552 338014
rect 362868 336728 362920 336734
rect 362868 336670 362920 336676
rect 363512 336728 363564 336734
rect 363512 336670 363564 336676
rect 363604 336524 363656 336530
rect 363604 336466 363656 336472
rect 362868 330540 362920 330546
rect 362868 330482 362920 330488
rect 362776 4820 362828 4826
rect 362776 4762 362828 4768
rect 361120 3528 361172 3534
rect 361120 3470 361172 3476
rect 361488 3528 361540 3534
rect 361488 3470 361540 3476
rect 361132 480 361160 3470
rect 362880 3466 362908 330482
rect 363616 5574 363644 336466
rect 363892 336190 363920 338014
rect 363880 336184 363932 336190
rect 363880 336126 363932 336132
rect 364168 7138 364196 338014
rect 364248 336728 364300 336734
rect 364248 336670 364300 336676
rect 364156 7132 364208 7138
rect 364156 7074 364208 7080
rect 363604 5568 363656 5574
rect 363604 5510 363656 5516
rect 363512 3732 363564 3738
rect 363512 3674 363564 3680
rect 362316 3460 362368 3466
rect 362316 3402 362368 3408
rect 362868 3460 362920 3466
rect 362868 3402 362920 3408
rect 362328 480 362356 3402
rect 363524 480 363552 3674
rect 364260 2854 364288 336670
rect 364628 335918 364656 338014
rect 364616 335912 364668 335918
rect 364616 335854 364668 335860
rect 364996 335578 365024 338014
rect 364984 335572 365036 335578
rect 364984 335514 365036 335520
rect 365364 335354 365392 338014
rect 365364 335326 365576 335354
rect 365548 7206 365576 335326
rect 365536 7200 365588 7206
rect 365536 7142 365588 7148
rect 364616 3188 364668 3194
rect 364616 3130 364668 3136
rect 364248 2848 364300 2854
rect 364248 2790 364300 2796
rect 364628 480 364656 3130
rect 365640 2922 365668 338014
rect 366100 335646 366128 338014
rect 366468 335850 366496 338014
rect 366456 335844 366508 335850
rect 366456 335786 366508 335792
rect 366836 335782 366864 338014
rect 366928 338014 366988 338042
rect 367264 338014 367508 338042
rect 367632 338014 367876 338042
rect 368000 338014 368244 338042
rect 366824 335776 366876 335782
rect 366824 335718 366876 335724
rect 366088 335640 366140 335646
rect 366088 335582 366140 335588
rect 366928 335510 366956 338014
rect 367376 336320 367428 336326
rect 367376 336262 367428 336268
rect 367008 335844 367060 335850
rect 367008 335786 367060 335792
rect 366916 335504 366968 335510
rect 366916 335446 366968 335452
rect 367020 7274 367048 335786
rect 367388 335354 367416 336262
rect 367480 335850 367508 338014
rect 367848 336462 367876 338014
rect 367836 336456 367888 336462
rect 367836 336398 367888 336404
rect 368216 336326 368244 338014
rect 368354 337770 368382 338028
rect 368736 338014 368980 338042
rect 369104 338014 369348 338042
rect 369472 338014 369716 338042
rect 368354 337742 368428 337770
rect 368204 336320 368256 336326
rect 368204 336262 368256 336268
rect 367468 335844 367520 335850
rect 367468 335786 367520 335792
rect 368296 335844 368348 335850
rect 368296 335786 368348 335792
rect 367388 335326 367508 335354
rect 367480 16574 367508 335326
rect 367480 16546 367784 16574
rect 367008 7268 367060 7274
rect 367008 7210 367060 7216
rect 367008 5568 367060 5574
rect 367008 5510 367060 5516
rect 365812 3256 365864 3262
rect 365812 3198 365864 3204
rect 365628 2916 365680 2922
rect 365628 2858 365680 2864
rect 365824 480 365852 3198
rect 367020 480 367048 5510
rect 367756 490 367784 16546
rect 368308 7342 368336 335786
rect 368400 7410 368428 337742
rect 368952 335714 368980 338014
rect 369320 335986 369348 338014
rect 369308 335980 369360 335986
rect 369308 335922 369360 335928
rect 368940 335708 368992 335714
rect 368940 335650 368992 335656
rect 369688 7478 369716 338014
rect 369780 338014 369840 338042
rect 370208 338014 370452 338042
rect 370576 338014 370820 338042
rect 370944 338014 371188 338042
rect 371312 338014 371556 338042
rect 371680 338014 371924 338042
rect 372048 338014 372292 338042
rect 369780 336666 369808 338014
rect 370424 336734 370452 338014
rect 370412 336728 370464 336734
rect 370412 336670 370464 336676
rect 369768 336660 369820 336666
rect 369768 336602 369820 336608
rect 370504 336388 370556 336394
rect 370504 336330 370556 336336
rect 369768 335708 369820 335714
rect 369768 335650 369820 335656
rect 369676 7472 369728 7478
rect 369676 7414 369728 7420
rect 368388 7404 368440 7410
rect 368388 7346 368440 7352
rect 368296 7336 368348 7342
rect 368296 7278 368348 7284
rect 369400 3324 369452 3330
rect 369400 3266 369452 3272
rect 368032 598 368244 626
rect 368032 490 368060 598
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 462 368060 490
rect 368216 480 368244 598
rect 369412 480 369440 3266
rect 369780 2990 369808 335650
rect 370516 6186 370544 336330
rect 370792 335354 370820 338014
rect 370792 335326 371096 335354
rect 370596 9036 370648 9042
rect 370596 8978 370648 8984
rect 370504 6180 370556 6186
rect 370504 6122 370556 6128
rect 369768 2984 369820 2990
rect 369768 2926 369820 2932
rect 370608 480 370636 8978
rect 371068 7546 371096 335326
rect 371056 7540 371108 7546
rect 371056 7482 371108 7488
rect 371160 3058 371188 338014
rect 371528 334490 371556 338014
rect 371792 336252 371844 336258
rect 371792 336194 371844 336200
rect 371804 335354 371832 336194
rect 371896 335578 371924 338014
rect 372264 336598 372292 338014
rect 372402 337770 372430 338028
rect 372784 338014 373028 338042
rect 373152 338014 373396 338042
rect 373520 338014 373764 338042
rect 372402 337742 372476 337770
rect 372252 336592 372304 336598
rect 372252 336534 372304 336540
rect 371884 335572 371936 335578
rect 371884 335514 371936 335520
rect 372344 335572 372396 335578
rect 372344 335514 372396 335520
rect 371804 335326 371924 335354
rect 371516 334484 371568 334490
rect 371516 334426 371568 334432
rect 371896 6254 371924 335326
rect 372356 8294 372384 335514
rect 372448 9042 372476 337742
rect 373000 335918 373028 338014
rect 373368 336530 373396 338014
rect 373356 336524 373408 336530
rect 373356 336466 373408 336472
rect 373736 336258 373764 338014
rect 373828 338014 373888 338042
rect 374256 338014 374500 338042
rect 374624 338014 374868 338042
rect 373724 336252 373776 336258
rect 373724 336194 373776 336200
rect 372988 335912 373040 335918
rect 372988 335854 373040 335860
rect 373828 333878 373856 338014
rect 373908 336524 373960 336530
rect 373908 336466 373960 336472
rect 373816 333872 373868 333878
rect 373816 333814 373868 333820
rect 372436 9036 372488 9042
rect 372436 8978 372488 8984
rect 372344 8288 372396 8294
rect 372344 8230 372396 8236
rect 371884 6248 371936 6254
rect 371884 6190 371936 6196
rect 372896 4072 372948 4078
rect 372896 4014 372948 4020
rect 371700 3392 371752 3398
rect 371700 3334 371752 3340
rect 371148 3052 371200 3058
rect 371148 2994 371200 3000
rect 371712 480 371740 3334
rect 372908 480 372936 4014
rect 373920 3126 373948 336466
rect 374472 336394 374500 338014
rect 374840 336530 374868 338014
rect 374978 337770 375006 338028
rect 375116 338014 375360 338042
rect 375728 338014 375972 338042
rect 376096 338014 376248 338042
rect 376464 338014 376616 338042
rect 376832 338014 377076 338042
rect 377200 338014 377444 338042
rect 377568 338014 377812 338042
rect 374978 337742 375052 337770
rect 374828 336524 374880 336530
rect 374828 336466 374880 336472
rect 374460 336388 374512 336394
rect 374460 336330 374512 336336
rect 374276 336252 374328 336258
rect 374276 336194 374328 336200
rect 374288 334558 374316 336194
rect 374644 335912 374696 335918
rect 374644 335854 374696 335860
rect 374276 334552 374328 334558
rect 374276 334494 374328 334500
rect 374656 333946 374684 335854
rect 374644 333940 374696 333946
rect 374644 333882 374696 333888
rect 375024 333810 375052 337742
rect 375012 333804 375064 333810
rect 375012 333746 375064 333752
rect 374092 4480 374144 4486
rect 374092 4422 374144 4428
rect 373908 3120 373960 3126
rect 373908 3062 373960 3068
rect 374104 480 374132 4422
rect 375116 3194 375144 338014
rect 375944 336530 375972 338014
rect 375196 336524 375248 336530
rect 375196 336466 375248 336472
rect 375932 336524 375984 336530
rect 375932 336466 375984 336472
rect 375208 5710 375236 336466
rect 375472 336116 375524 336122
rect 375472 336058 375524 336064
rect 375484 16574 375512 336058
rect 376220 332382 376248 338014
rect 376588 336258 376616 338014
rect 377048 336530 377076 338014
rect 376668 336524 376720 336530
rect 376668 336466 376720 336472
rect 377036 336524 377088 336530
rect 377036 336466 377088 336472
rect 376576 336252 376628 336258
rect 376576 336194 376628 336200
rect 376208 332376 376260 332382
rect 376208 332318 376260 332324
rect 375484 16546 376064 16574
rect 375196 5704 375248 5710
rect 375196 5646 375248 5652
rect 375288 4140 375340 4146
rect 375288 4082 375340 4088
rect 375104 3188 375156 3194
rect 375104 3130 375156 3136
rect 375300 480 375328 4082
rect 376036 490 376064 16546
rect 376680 5778 376708 336466
rect 377416 333742 377444 338014
rect 377404 333736 377456 333742
rect 377404 333678 377456 333684
rect 376668 5772 376720 5778
rect 376668 5714 376720 5720
rect 377680 4548 377732 4554
rect 377680 4490 377732 4496
rect 376312 598 376524 626
rect 376312 490 376340 598
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 462 376340 490
rect 376496 480 376524 598
rect 377692 480 377720 4490
rect 377784 3262 377812 338014
rect 377922 337770 377950 338028
rect 378304 338014 378548 338042
rect 378672 338014 378916 338042
rect 379040 338014 379192 338042
rect 379316 338014 379468 338042
rect 379684 338014 379928 338042
rect 380052 338014 380296 338042
rect 380420 338014 380572 338042
rect 377922 337742 377996 337770
rect 377864 336524 377916 336530
rect 377864 336466 377916 336472
rect 377876 5846 377904 336466
rect 377968 5914 377996 337742
rect 378520 332314 378548 338014
rect 378888 336394 378916 338014
rect 378876 336388 378928 336394
rect 378876 336330 378928 336336
rect 378508 332308 378560 332314
rect 378508 332250 378560 332256
rect 379164 325694 379192 338014
rect 379440 332246 379468 338014
rect 379900 336462 379928 338014
rect 380268 336530 380296 338014
rect 380256 336524 380308 336530
rect 380256 336466 380308 336472
rect 379888 336456 379940 336462
rect 379888 336398 379940 336404
rect 380544 333674 380572 338014
rect 380774 337770 380802 338028
rect 381156 338014 381400 338042
rect 381524 338014 381768 338042
rect 381892 338014 382136 338042
rect 380774 337742 380848 337770
rect 380716 336524 380768 336530
rect 380716 336466 380768 336472
rect 380624 336456 380676 336462
rect 380624 336398 380676 336404
rect 380532 333668 380584 333674
rect 380532 333610 380584 333616
rect 379428 332240 379480 332246
rect 379428 332182 379480 332188
rect 379164 325666 379468 325694
rect 378876 6248 378928 6254
rect 378876 6190 378928 6196
rect 377956 5908 378008 5914
rect 377956 5850 378008 5856
rect 377864 5840 377916 5846
rect 377864 5782 377916 5788
rect 377772 3256 377824 3262
rect 377772 3198 377824 3204
rect 378888 480 378916 6190
rect 379440 5982 379468 325666
rect 379428 5976 379480 5982
rect 379428 5918 379480 5924
rect 379980 4004 380032 4010
rect 379980 3946 380032 3952
rect 379992 480 380020 3946
rect 380636 3330 380664 336398
rect 380728 6050 380756 336466
rect 380820 336258 380848 337742
rect 380808 336252 380860 336258
rect 380808 336194 380860 336200
rect 381372 330546 381400 338014
rect 381740 336326 381768 338014
rect 382004 336524 382056 336530
rect 382004 336466 382056 336472
rect 381728 336320 381780 336326
rect 381728 336262 381780 336268
rect 381360 330540 381412 330546
rect 381360 330482 381412 330488
rect 382016 6798 382044 336466
rect 382108 335354 382136 338014
rect 382200 338014 382260 338042
rect 382628 338014 382872 338042
rect 382996 338014 383240 338042
rect 383364 338014 383516 338042
rect 383732 338014 383976 338042
rect 384100 338014 384344 338042
rect 384468 338014 384712 338042
rect 382200 336530 382228 338014
rect 382188 336524 382240 336530
rect 382188 336466 382240 336472
rect 382464 336048 382516 336054
rect 382464 335990 382516 335996
rect 382108 335326 382228 335354
rect 382096 330540 382148 330546
rect 382096 330482 382148 330488
rect 382004 6792 382056 6798
rect 382004 6734 382056 6740
rect 382108 6118 382136 330482
rect 382096 6112 382148 6118
rect 382096 6054 382148 6060
rect 380716 6044 380768 6050
rect 380716 5986 380768 5992
rect 381176 4616 381228 4622
rect 381176 4558 381228 4564
rect 380624 3324 380676 3330
rect 380624 3266 380676 3272
rect 381188 480 381216 4558
rect 382200 3398 382228 335326
rect 382372 8968 382424 8974
rect 382372 8910 382424 8916
rect 382188 3392 382240 3398
rect 382188 3334 382240 3340
rect 382384 480 382412 8910
rect 382476 6914 382504 335990
rect 382844 332178 382872 338014
rect 383212 336122 383240 338014
rect 383488 336190 383516 338014
rect 383476 336184 383528 336190
rect 383476 336126 383528 336132
rect 382924 336116 382976 336122
rect 382924 336058 382976 336064
rect 383200 336116 383252 336122
rect 383200 336058 383252 336064
rect 382832 332172 382884 332178
rect 382832 332114 382884 332120
rect 382936 8974 382964 336058
rect 383948 336054 383976 338014
rect 383936 336048 383988 336054
rect 383936 335990 383988 335996
rect 384316 335238 384344 338014
rect 384684 336705 384712 338014
rect 384776 338014 384836 338042
rect 385204 338014 385356 338042
rect 385572 338014 385816 338042
rect 385940 338014 386184 338042
rect 384670 336696 384726 336705
rect 384670 336631 384726 336640
rect 384304 335232 384356 335238
rect 384304 335174 384356 335180
rect 382924 8968 382976 8974
rect 382924 8910 382976 8916
rect 382476 6886 383608 6914
rect 383580 480 383608 6886
rect 384776 6662 384804 338014
rect 384856 336048 384908 336054
rect 384856 335990 384908 335996
rect 384868 6730 384896 335990
rect 385328 332110 385356 338014
rect 385788 336161 385816 338014
rect 385774 336152 385830 336161
rect 385774 336087 385830 336096
rect 385316 332104 385368 332110
rect 385316 332046 385368 332052
rect 386156 325694 386184 338014
rect 386294 337770 386322 338028
rect 386676 338014 386920 338042
rect 387044 338014 387288 338042
rect 387412 338014 387656 338042
rect 386294 337742 386368 337770
rect 386340 332042 386368 337742
rect 386892 336569 386920 338014
rect 386878 336560 386934 336569
rect 386878 336495 386934 336504
rect 387260 336054 387288 338014
rect 387248 336048 387300 336054
rect 387248 335990 387300 335996
rect 387628 333606 387656 338014
rect 387720 338014 387780 338042
rect 388148 338014 388392 338042
rect 388516 338014 388760 338042
rect 387720 336297 387748 338014
rect 387706 336288 387762 336297
rect 387706 336223 387762 336232
rect 388364 336054 388392 338014
rect 387708 336048 387760 336054
rect 387708 335990 387760 335996
rect 388352 336048 388404 336054
rect 388352 335990 388404 335996
rect 387616 333600 387668 333606
rect 387616 333542 387668 333548
rect 386328 332036 386380 332042
rect 386328 331978 386380 331984
rect 386156 325666 386368 325694
rect 384856 6724 384908 6730
rect 384856 6666 384908 6672
rect 384764 6656 384816 6662
rect 384764 6598 384816 6604
rect 386340 6594 386368 325666
rect 386328 6588 386380 6594
rect 386328 6530 386380 6536
rect 387720 6526 387748 335990
rect 388444 335368 388496 335374
rect 388444 335310 388496 335316
rect 387708 6520 387760 6526
rect 387708 6462 387760 6468
rect 385960 6180 386012 6186
rect 385960 6122 386012 6128
rect 384764 4684 384816 4690
rect 384764 4626 384816 4632
rect 384776 480 384804 4626
rect 385972 480 386000 6122
rect 388260 4752 388312 4758
rect 388260 4694 388312 4700
rect 387156 3936 387208 3942
rect 387156 3878 387208 3884
rect 387168 480 387196 3878
rect 388272 480 388300 4694
rect 388456 4214 388484 335310
rect 388732 331974 388760 338014
rect 388824 338014 388884 338042
rect 389252 338014 389496 338042
rect 389620 338014 389864 338042
rect 389988 338014 390140 338042
rect 388824 335374 388852 338014
rect 388994 336696 389050 336705
rect 388994 336631 389050 336640
rect 388812 335368 388864 335374
rect 388812 335310 388864 335316
rect 389008 335306 389036 336631
rect 389468 336054 389496 338014
rect 389088 336048 389140 336054
rect 389088 335990 389140 335996
rect 389456 336048 389508 336054
rect 389456 335990 389508 335996
rect 388996 335300 389048 335306
rect 388996 335242 389048 335248
rect 388720 331968 388772 331974
rect 388720 331910 388772 331916
rect 389100 6458 389128 335990
rect 389836 330818 389864 338014
rect 390112 335102 390140 338014
rect 390342 337770 390370 338028
rect 390724 338014 390968 338042
rect 391092 338014 391244 338042
rect 391368 338014 391612 338042
rect 391736 338014 391888 338042
rect 392104 338014 392348 338042
rect 392472 338014 392716 338042
rect 390342 337742 390416 337770
rect 390192 336048 390244 336054
rect 390192 335990 390244 335996
rect 390100 335096 390152 335102
rect 390100 335038 390152 335044
rect 389824 330812 389876 330818
rect 389824 330754 389876 330760
rect 389088 6452 389140 6458
rect 389088 6394 389140 6400
rect 390204 6390 390232 335990
rect 390192 6384 390244 6390
rect 390192 6326 390244 6332
rect 390388 6322 390416 337742
rect 390940 333538 390968 338014
rect 391216 336025 391244 338014
rect 391202 336016 391258 336025
rect 391202 335951 391258 335960
rect 391584 335354 391612 338014
rect 391584 335326 391704 335354
rect 390928 333532 390980 333538
rect 390928 333474 390980 333480
rect 390376 6316 390428 6322
rect 390376 6258 390428 6264
rect 391676 6254 391704 335326
rect 391860 331906 391888 338014
rect 391938 336560 391994 336569
rect 391938 336495 391994 336504
rect 391952 335170 391980 336495
rect 391940 335164 391992 335170
rect 391940 335106 391992 335112
rect 392320 335034 392348 338014
rect 392688 336054 392716 338014
rect 392826 337770 392854 338028
rect 392964 338014 393208 338042
rect 393576 338014 393820 338042
rect 393944 338014 394188 338042
rect 394312 338014 394464 338042
rect 392826 337742 392900 337770
rect 392676 336048 392728 336054
rect 392676 335990 392728 335996
rect 392308 335028 392360 335034
rect 392308 334970 392360 334976
rect 391848 331900 391900 331906
rect 391848 331842 391900 331848
rect 392872 330750 392900 337742
rect 392860 330744 392912 330750
rect 392860 330686 392912 330692
rect 392584 10328 392636 10334
rect 392584 10270 392636 10276
rect 391664 6248 391716 6254
rect 391664 6190 391716 6196
rect 391848 5500 391900 5506
rect 391848 5442 391900 5448
rect 388444 4208 388496 4214
rect 388444 4150 388496 4156
rect 389456 4208 389508 4214
rect 389456 4150 389508 4156
rect 389468 480 389496 4150
rect 390652 3868 390704 3874
rect 390652 3810 390704 3816
rect 390664 480 390692 3810
rect 391860 480 391888 5442
rect 392596 490 392624 10270
rect 392964 4282 392992 338014
rect 393136 336048 393188 336054
rect 393136 335990 393188 335996
rect 393148 6186 393176 335990
rect 393792 334966 393820 338014
rect 393780 334960 393832 334966
rect 393780 334902 393832 334908
rect 394160 330682 394188 338014
rect 394148 330676 394200 330682
rect 394148 330618 394200 330624
rect 393136 6180 393188 6186
rect 393136 6122 393188 6128
rect 394436 4350 394464 338014
rect 394620 338014 394680 338042
rect 395048 338014 395200 338042
rect 395416 338014 395660 338042
rect 395784 338014 395936 338042
rect 396152 338014 396396 338042
rect 396520 338014 396764 338042
rect 396888 338014 397132 338042
rect 397256 338014 397408 338042
rect 397624 338014 397868 338042
rect 397992 338014 398236 338042
rect 398360 338014 398512 338042
rect 394620 333470 394648 338014
rect 394608 333464 394660 333470
rect 394608 333406 394660 333412
rect 395172 330614 395200 338014
rect 395344 336048 395396 336054
rect 395344 335990 395396 335996
rect 395160 330608 395212 330614
rect 395160 330550 395212 330556
rect 395252 5432 395304 5438
rect 395252 5374 395304 5380
rect 394424 4344 394476 4350
rect 394424 4286 394476 4292
rect 392952 4276 393004 4282
rect 392952 4218 393004 4224
rect 394240 3800 394292 3806
rect 394240 3742 394292 3748
rect 392872 598 393084 626
rect 392872 490 392900 598
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 462 392900 490
rect 393056 480 393084 598
rect 394252 480 394280 3742
rect 395264 2802 395292 5374
rect 395356 4214 395384 335990
rect 395632 335354 395660 338014
rect 395632 335326 395844 335354
rect 395816 4418 395844 335326
rect 395908 334898 395936 338014
rect 395896 334892 395948 334898
rect 395896 334834 395948 334840
rect 396368 330546 396396 338014
rect 396356 330540 396408 330546
rect 396356 330482 396408 330488
rect 396736 325694 396764 338014
rect 397104 334762 397132 338014
rect 397092 334756 397144 334762
rect 397092 334698 397144 334704
rect 397380 329186 397408 338014
rect 397840 336054 397868 338014
rect 397828 336048 397880 336054
rect 397828 335990 397880 335996
rect 398208 334830 398236 338014
rect 398196 334824 398248 334830
rect 398196 334766 398248 334772
rect 398484 334694 398512 338014
rect 398668 338014 398728 338042
rect 399096 338014 399340 338042
rect 399464 338014 399708 338042
rect 398564 336048 398616 336054
rect 398564 335990 398616 335996
rect 398472 334688 398524 334694
rect 398472 334630 398524 334636
rect 397368 329180 397420 329186
rect 397368 329122 397420 329128
rect 396736 325666 397132 325694
rect 397104 4486 397132 325666
rect 398576 4554 398604 335990
rect 398668 4622 398696 338014
rect 399312 333402 399340 338014
rect 399300 333396 399352 333402
rect 399300 333338 399352 333344
rect 399680 330886 399708 338014
rect 399818 337770 399846 338028
rect 400140 338014 400200 338042
rect 400568 338014 400812 338042
rect 400936 338014 401180 338042
rect 401304 338014 401548 338042
rect 401672 338014 401916 338042
rect 402040 338014 402284 338042
rect 402408 338014 402560 338042
rect 399818 337742 399892 337770
rect 399668 330880 399720 330886
rect 399668 330822 399720 330828
rect 398932 5296 398984 5302
rect 398932 5238 398984 5244
rect 398656 4616 398708 4622
rect 398656 4558 398708 4564
rect 398564 4548 398616 4554
rect 398564 4490 398616 4496
rect 397092 4480 397144 4486
rect 397092 4422 397144 4428
rect 395804 4412 395856 4418
rect 395804 4354 395856 4360
rect 395344 4208 395396 4214
rect 395344 4150 395396 4156
rect 396540 4208 396592 4214
rect 396540 4150 396592 4156
rect 395264 2774 395384 2802
rect 395356 480 395384 2774
rect 396552 480 396580 4150
rect 397736 3732 397788 3738
rect 397736 3674 397788 3680
rect 397748 480 397776 3674
rect 398944 480 398972 5238
rect 399864 4690 399892 337742
rect 400140 333334 400168 338014
rect 400128 333328 400180 333334
rect 400128 333270 400180 333276
rect 400784 329118 400812 338014
rect 401152 335354 401180 338014
rect 401152 335326 401364 335354
rect 400772 329112 400824 329118
rect 400772 329054 400824 329060
rect 400128 5364 400180 5370
rect 400128 5306 400180 5312
rect 399852 4684 399904 4690
rect 399852 4626 399904 4632
rect 400140 480 400168 5306
rect 401336 4758 401364 335326
rect 401520 333266 401548 338014
rect 401888 335442 401916 338014
rect 402256 336054 402284 338014
rect 402244 336048 402296 336054
rect 402244 335990 402296 335996
rect 401876 335436 401928 335442
rect 401876 335378 401928 335384
rect 402532 334626 402560 338014
rect 402762 337770 402790 338028
rect 403144 338014 403296 338042
rect 403420 338014 403664 338042
rect 403788 338014 404032 338042
rect 402762 337742 402836 337770
rect 402704 336048 402756 336054
rect 402704 335990 402756 335996
rect 402612 335436 402664 335442
rect 402612 335378 402664 335384
rect 402520 334620 402572 334626
rect 402520 334562 402572 334568
rect 401508 333260 401560 333266
rect 401508 333202 401560 333208
rect 402520 5228 402572 5234
rect 402520 5170 402572 5176
rect 401324 4752 401376 4758
rect 401324 4694 401376 4700
rect 401324 3664 401376 3670
rect 401324 3606 401376 3612
rect 401336 480 401364 3606
rect 402532 480 402560 5170
rect 402624 4146 402652 335378
rect 402716 5506 402744 335990
rect 402704 5500 402756 5506
rect 402704 5442 402756 5448
rect 402612 4140 402664 4146
rect 402612 4082 402664 4088
rect 402808 4078 402836 337742
rect 403268 335374 403296 338014
rect 403256 335368 403308 335374
rect 403256 335310 403308 335316
rect 403636 325694 403664 338014
rect 404004 335442 404032 338014
rect 404096 338014 404156 338042
rect 404524 338014 404768 338042
rect 404892 338014 405136 338042
rect 405260 338014 405412 338042
rect 403992 335436 404044 335442
rect 403992 335378 404044 335384
rect 403636 325666 404032 325694
rect 404004 8226 404032 325666
rect 403992 8220 404044 8226
rect 403992 8162 404044 8168
rect 404096 5370 404124 338014
rect 404740 335442 404768 338014
rect 404268 335436 404320 335442
rect 404268 335378 404320 335384
rect 404728 335436 404780 335442
rect 404728 335378 404780 335384
rect 404176 335368 404228 335374
rect 404176 335310 404228 335316
rect 404188 5438 404216 335310
rect 404176 5432 404228 5438
rect 404176 5374 404228 5380
rect 404084 5364 404136 5370
rect 404084 5306 404136 5312
rect 403624 5160 403676 5166
rect 403624 5102 403676 5108
rect 402796 4072 402848 4078
rect 402796 4014 402848 4020
rect 403636 480 403664 5102
rect 404280 4010 404308 335378
rect 405108 335374 405136 338014
rect 405384 335442 405412 338014
rect 405476 338014 405628 338042
rect 405996 338014 406240 338042
rect 406364 338014 406608 338042
rect 405280 335436 405332 335442
rect 405280 335378 405332 335384
rect 405372 335436 405424 335442
rect 405372 335378 405424 335384
rect 405096 335368 405148 335374
rect 405096 335310 405148 335316
rect 405292 325694 405320 335378
rect 405292 325666 405412 325694
rect 405384 8158 405412 325666
rect 405372 8152 405424 8158
rect 405372 8094 405424 8100
rect 405476 8090 405504 338014
rect 405556 335436 405608 335442
rect 405556 335378 405608 335384
rect 405464 8084 405516 8090
rect 405464 8026 405516 8032
rect 405568 5302 405596 335378
rect 406212 335374 406240 338014
rect 406580 335442 406608 338014
rect 406718 337770 406746 338028
rect 406948 338014 407100 338042
rect 407468 338014 407712 338042
rect 407836 338014 408080 338042
rect 408204 338014 408448 338042
rect 408572 338014 408816 338042
rect 408940 338014 409184 338042
rect 409308 338014 409552 338042
rect 406718 337742 406792 337770
rect 406568 335436 406620 335442
rect 406568 335378 406620 335384
rect 405648 335368 405700 335374
rect 405648 335310 405700 335316
rect 406200 335368 406252 335374
rect 406200 335310 406252 335316
rect 405556 5296 405608 5302
rect 405556 5238 405608 5244
rect 404268 4004 404320 4010
rect 404268 3946 404320 3952
rect 405660 3942 405688 335310
rect 406764 8022 406792 337742
rect 406844 335436 406896 335442
rect 406844 335378 406896 335384
rect 406752 8016 406804 8022
rect 406752 7958 406804 7964
rect 406856 5234 406884 335378
rect 406844 5228 406896 5234
rect 406844 5170 406896 5176
rect 406016 5092 406068 5098
rect 406016 5034 406068 5040
rect 405648 3936 405700 3942
rect 405648 3878 405700 3884
rect 404820 3596 404872 3602
rect 404820 3538 404872 3544
rect 404832 480 404860 3538
rect 406028 480 406056 5034
rect 406948 3806 406976 338014
rect 407684 335442 407712 338014
rect 407672 335436 407724 335442
rect 407672 335378 407724 335384
rect 407028 335368 407080 335374
rect 408052 335354 408080 338014
rect 408316 335436 408368 335442
rect 408316 335378 408368 335384
rect 408052 335326 408264 335354
rect 407028 335310 407080 335316
rect 407040 3874 407068 335310
rect 408236 7954 408264 335326
rect 408224 7948 408276 7954
rect 408224 7890 408276 7896
rect 408328 5166 408356 335378
rect 408316 5160 408368 5166
rect 408316 5102 408368 5108
rect 407212 5024 407264 5030
rect 407212 4966 407264 4972
rect 407028 3868 407080 3874
rect 407028 3810 407080 3816
rect 406936 3800 406988 3806
rect 406936 3742 406988 3748
rect 407224 480 407252 4966
rect 408420 3738 408448 338014
rect 408788 335374 408816 338014
rect 408776 335368 408828 335374
rect 408776 335310 408828 335316
rect 409156 325694 409184 338014
rect 409524 335442 409552 338014
rect 409662 337770 409690 338028
rect 410044 338014 410288 338042
rect 410412 338014 410656 338042
rect 409662 337742 409736 337770
rect 409512 335436 409564 335442
rect 409512 335378 409564 335384
rect 409604 335368 409656 335374
rect 409604 335310 409656 335316
rect 409156 325666 409552 325694
rect 409524 7886 409552 325666
rect 409512 7880 409564 7886
rect 409512 7822 409564 7828
rect 409616 5098 409644 335310
rect 409604 5092 409656 5098
rect 409604 5034 409656 5040
rect 409708 5030 409736 337742
rect 409788 335436 409840 335442
rect 409788 335378 409840 335384
rect 409696 5024 409748 5030
rect 409696 4966 409748 4972
rect 409604 4888 409656 4894
rect 409604 4830 409656 4836
rect 408408 3732 408460 3738
rect 408408 3674 408460 3680
rect 408408 3528 408460 3534
rect 408408 3470 408460 3476
rect 408420 480 408448 3470
rect 409616 480 409644 4830
rect 409800 3670 409828 335378
rect 410260 335374 410288 338014
rect 410248 335368 410300 335374
rect 410248 335310 410300 335316
rect 410628 331158 410656 338014
rect 410720 338014 410780 338042
rect 410904 338014 411148 338042
rect 411516 338014 411760 338042
rect 411884 338014 412128 338042
rect 410720 335442 410748 338014
rect 410708 335436 410760 335442
rect 410708 335378 410760 335384
rect 410616 331152 410668 331158
rect 410616 331094 410668 331100
rect 410904 7750 410932 338014
rect 411076 335436 411128 335442
rect 411076 335378 411128 335384
rect 410984 335368 411036 335374
rect 410984 335310 411036 335316
rect 410996 7818 411024 335310
rect 410984 7812 411036 7818
rect 410984 7754 411036 7760
rect 410892 7744 410944 7750
rect 410892 7686 410944 7692
rect 411088 4962 411116 335378
rect 411732 335374 411760 338014
rect 412100 335442 412128 338014
rect 412238 337770 412266 338028
rect 412560 338014 412620 338042
rect 412988 338014 413232 338042
rect 413356 338014 413600 338042
rect 413724 338014 413968 338042
rect 414092 338014 414336 338042
rect 414460 338014 414704 338042
rect 412238 337742 412312 337770
rect 412088 335436 412140 335442
rect 412088 335378 412140 335384
rect 411720 335368 411772 335374
rect 411720 335310 411772 335316
rect 411168 331152 411220 331158
rect 411168 331094 411220 331100
rect 410800 4956 410852 4962
rect 410800 4898 410852 4904
rect 411076 4956 411128 4962
rect 411076 4898 411128 4904
rect 409788 3664 409840 3670
rect 409788 3606 409840 3612
rect 410812 480 410840 4898
rect 411180 3602 411208 331094
rect 412284 7682 412312 337742
rect 412364 335436 412416 335442
rect 412364 335378 412416 335384
rect 412272 7676 412324 7682
rect 412272 7618 412324 7624
rect 412376 4894 412404 335378
rect 412456 335368 412508 335374
rect 412456 335310 412508 335316
rect 412364 4888 412416 4894
rect 412364 4830 412416 4836
rect 411168 3596 411220 3602
rect 411168 3538 411220 3544
rect 412468 3534 412496 335310
rect 412456 3528 412508 3534
rect 412456 3470 412508 3476
rect 412560 3466 412588 338014
rect 413204 335714 413232 338014
rect 413192 335708 413244 335714
rect 413192 335650 413244 335656
rect 413572 335354 413600 338014
rect 413836 335708 413888 335714
rect 413836 335650 413888 335656
rect 413572 335326 413784 335354
rect 413756 7614 413784 335326
rect 413744 7608 413796 7614
rect 413744 7550 413796 7556
rect 413848 4826 413876 335650
rect 413100 4820 413152 4826
rect 413100 4762 413152 4768
rect 413836 4820 413888 4826
rect 413836 4762 413888 4768
rect 411904 3460 411956 3466
rect 411904 3402 411956 3408
rect 412548 3460 412600 3466
rect 412548 3402 412600 3408
rect 411916 480 411944 3402
rect 413112 480 413140 4762
rect 413940 3777 413968 338014
rect 414308 330478 414336 338014
rect 414676 335646 414704 338014
rect 414768 338014 414828 338042
rect 414768 335714 414796 338014
rect 414756 335708 414808 335714
rect 414756 335650 414808 335656
rect 414664 335640 414716 335646
rect 414664 335582 414716 335588
rect 414296 330472 414348 330478
rect 414296 330414 414348 330420
rect 414952 20670 414980 457286
rect 417424 457224 417476 457230
rect 417424 457166 417476 457172
rect 417436 353258 417464 457166
rect 418816 405686 418844 458662
rect 428464 458652 428516 458658
rect 428464 458594 428516 458600
rect 421656 458516 421708 458522
rect 421656 458458 421708 458464
rect 418804 405680 418856 405686
rect 418804 405622 418856 405628
rect 417424 353252 417476 353258
rect 417424 353194 417476 353200
rect 417422 336288 417478 336297
rect 417422 336223 417478 336232
rect 415308 335708 415360 335714
rect 415308 335650 415360 335656
rect 415216 335640 415268 335646
rect 415216 335582 415268 335588
rect 415124 330472 415176 330478
rect 415124 330414 415176 330420
rect 414940 20664 414992 20670
rect 414940 20606 414992 20612
rect 414296 7064 414348 7070
rect 414296 7006 414348 7012
rect 413926 3768 413982 3777
rect 413926 3703 413982 3712
rect 414308 480 414336 7006
rect 415136 3505 415164 330414
rect 415228 3641 415256 335582
rect 415214 3632 415270 3641
rect 415214 3567 415270 3576
rect 415122 3496 415178 3505
rect 415122 3431 415178 3440
rect 415320 3369 415348 335650
rect 417436 8974 417464 336223
rect 417516 335572 417568 335578
rect 417516 335514 417568 335520
rect 417528 9654 417556 335514
rect 418804 335504 418856 335510
rect 418804 335446 418856 335452
rect 418160 335436 418212 335442
rect 418160 335378 418212 335384
rect 418172 16574 418200 335378
rect 418172 16546 418568 16574
rect 417516 9648 417568 9654
rect 417516 9590 417568 9596
rect 416688 8968 416740 8974
rect 416688 8910 416740 8916
rect 417424 8968 417476 8974
rect 417424 8910 417476 8916
rect 415306 3360 415362 3369
rect 415306 3295 415362 3304
rect 415492 2848 415544 2854
rect 415492 2790 415544 2796
rect 415504 480 415532 2790
rect 416700 480 416728 8910
rect 417884 7132 417936 7138
rect 417884 7074 417936 7080
rect 417896 480 417924 7074
rect 418540 490 418568 16546
rect 418816 9110 418844 335446
rect 421564 335368 421616 335374
rect 421564 335310 421616 335316
rect 420184 9648 420236 9654
rect 420184 9590 420236 9596
rect 418804 9104 418856 9110
rect 418804 9046 418856 9052
rect 418816 598 419028 626
rect 418816 490 418844 598
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418540 462 418844 490
rect 419000 480 419028 598
rect 420196 480 420224 9590
rect 421576 8362 421604 335310
rect 421668 325650 421696 458458
rect 425704 457156 425756 457162
rect 425704 457098 425756 457104
rect 425716 379506 425744 457098
rect 428476 431934 428504 458594
rect 429844 458380 429896 458386
rect 429844 458322 429896 458328
rect 428464 431928 428516 431934
rect 428464 431870 428516 431876
rect 425704 379500 425756 379506
rect 425704 379442 425756 379448
rect 429856 365702 429884 458322
rect 431224 456952 431276 456958
rect 431224 456894 431276 456900
rect 429844 365696 429896 365702
rect 429844 365638 429896 365644
rect 429200 335912 429252 335918
rect 429200 335854 429252 335860
rect 428464 335844 428516 335850
rect 428464 335786 428516 335792
rect 425060 335776 425112 335782
rect 425060 335718 425112 335724
rect 421656 325644 421708 325650
rect 421656 325586 421708 325592
rect 425072 16574 425100 335718
rect 425072 16546 425744 16574
rect 421564 8356 421616 8362
rect 421564 8298 421616 8304
rect 423772 8356 423824 8362
rect 423772 8298 423824 8304
rect 421380 7200 421432 7206
rect 421380 7142 421432 7148
rect 421392 480 421420 7142
rect 422576 2916 422628 2922
rect 422576 2858 422628 2864
rect 422588 480 422616 2858
rect 423784 480 423812 8298
rect 424968 7268 425020 7274
rect 424968 7210 425020 7216
rect 424980 480 425008 7210
rect 425716 490 425744 16546
rect 428476 11014 428504 335786
rect 428464 11008 428516 11014
rect 428464 10950 428516 10956
rect 427268 9104 427320 9110
rect 427268 9046 427320 9052
rect 425992 598 426204 626
rect 425992 490 426020 598
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 462 426020 490
rect 426176 480 426204 598
rect 427280 480 427308 9046
rect 428464 7336 428516 7342
rect 428464 7278 428516 7284
rect 428476 480 428504 7278
rect 429212 490 429240 335854
rect 431236 20670 431264 456894
rect 435364 336728 435416 336734
rect 435364 336670 435416 336676
rect 432604 335980 432656 335986
rect 432604 335922 432656 335928
rect 431224 20664 431276 20670
rect 431224 20606 431276 20612
rect 430856 11008 430908 11014
rect 430856 10950 430908 10956
rect 429488 598 429700 626
rect 429488 490 429516 598
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429212 462 429516 490
rect 429672 480 429700 598
rect 430868 480 430896 10950
rect 432616 7546 432644 335922
rect 435376 7546 435404 336670
rect 436100 336660 436152 336666
rect 436100 336602 436152 336608
rect 436112 16574 436140 336602
rect 443000 336592 443052 336598
rect 443000 336534 443052 336540
rect 440332 334484 440384 334490
rect 440332 334426 440384 334432
rect 436112 16546 436784 16574
rect 432604 7540 432656 7546
rect 432604 7482 432656 7488
rect 434444 7540 434496 7546
rect 434444 7482 434496 7488
rect 435364 7540 435416 7546
rect 435364 7482 435416 7488
rect 432052 7404 432104 7410
rect 432052 7346 432104 7352
rect 432064 480 432092 7346
rect 433248 2984 433300 2990
rect 433248 2926 433300 2932
rect 433260 480 433288 2926
rect 434456 480 434484 7482
rect 435548 7336 435600 7342
rect 435548 7278 435600 7284
rect 435560 480 435588 7278
rect 436756 480 436784 16546
rect 440344 11762 440372 334426
rect 443012 16574 443040 336534
rect 449900 336524 449952 336530
rect 449900 336466 449952 336472
rect 448520 334552 448572 334558
rect 448520 334494 448572 334500
rect 445760 333940 445812 333946
rect 445760 333882 445812 333888
rect 443012 16546 443408 16574
rect 440332 11756 440384 11762
rect 440332 11698 440384 11704
rect 441528 11756 441580 11762
rect 441528 11698 441580 11704
rect 437940 7540 437992 7546
rect 437940 7482 437992 7488
rect 437952 480 437980 7482
rect 439136 7404 439188 7410
rect 439136 7346 439188 7352
rect 439148 480 439176 7346
rect 440332 3052 440384 3058
rect 440332 2994 440384 3000
rect 440344 480 440372 2994
rect 441540 480 441568 11698
rect 442632 8288 442684 8294
rect 442632 8230 442684 8236
rect 442644 480 442672 8230
rect 443380 490 443408 16546
rect 445024 9036 445076 9042
rect 445024 8978 445076 8984
rect 443656 598 443868 626
rect 443656 490 443684 598
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 462 443684 490
rect 443840 480 443868 598
rect 445036 480 445064 8978
rect 445772 490 445800 333882
rect 448532 6914 448560 334494
rect 448612 333872 448664 333878
rect 448612 333814 448664 333820
rect 448624 11762 448652 333814
rect 449912 16574 449940 336466
rect 456800 336456 456852 336462
rect 456800 336398 456852 336404
rect 452660 333804 452712 333810
rect 452660 333746 452712 333752
rect 452672 16574 452700 333746
rect 449912 16546 450952 16574
rect 452672 16546 453344 16574
rect 448612 11756 448664 11762
rect 448612 11698 448664 11704
rect 449808 11756 449860 11762
rect 449808 11698 449860 11704
rect 448532 6886 448652 6914
rect 447416 3120 447468 3126
rect 447416 3062 447468 3068
rect 446048 598 446260 626
rect 446048 490 446076 598
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 462 446076 490
rect 446232 480 446260 598
rect 447428 480 447456 3062
rect 448624 480 448652 6886
rect 449820 480 449848 11698
rect 450924 480 450952 16546
rect 452108 5704 452160 5710
rect 452108 5646 452160 5652
rect 452120 480 452148 5646
rect 453316 480 453344 16546
rect 455696 5772 455748 5778
rect 455696 5714 455748 5720
rect 454500 3188 454552 3194
rect 454500 3130 454552 3136
rect 454512 480 454540 3130
rect 455708 480 455736 5714
rect 456812 3194 456840 336398
rect 465080 336388 465132 336394
rect 465080 336330 465132 336336
rect 459560 333736 459612 333742
rect 459560 333678 459612 333684
rect 456892 332376 456944 332382
rect 456892 332318 456944 332324
rect 456800 3188 456852 3194
rect 456800 3130 456852 3136
rect 456904 480 456932 332318
rect 459572 16574 459600 333678
rect 463700 332308 463752 332314
rect 463700 332250 463752 332256
rect 463712 16574 463740 332250
rect 465092 16574 465120 336330
rect 468484 336320 468536 336326
rect 468484 336262 468536 336268
rect 466460 332240 466512 332246
rect 466460 332182 466512 332188
rect 466472 16574 466500 332182
rect 459572 16546 459968 16574
rect 463712 16546 464016 16574
rect 465092 16546 465212 16574
rect 466472 16546 467512 16574
rect 459192 5840 459244 5846
rect 459192 5782 459244 5788
rect 458088 3188 458140 3194
rect 458088 3130 458140 3136
rect 458100 480 458128 3130
rect 459204 480 459232 5782
rect 459940 490 459968 16546
rect 462780 5908 462832 5914
rect 462780 5850 462832 5856
rect 461584 3256 461636 3262
rect 461584 3198 461636 3204
rect 460216 598 460428 626
rect 460216 490 460244 598
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 462 460244 490
rect 460400 480 460428 598
rect 461596 480 461624 3198
rect 462792 480 462820 5850
rect 463988 480 464016 16546
rect 465184 480 465212 16546
rect 466276 5976 466328 5982
rect 466276 5918 466328 5924
rect 466288 480 466316 5918
rect 467484 480 467512 16546
rect 468496 5982 468524 336262
rect 471980 336252 472032 336258
rect 471980 336194 472032 336200
rect 470600 333668 470652 333674
rect 470600 333610 470652 333616
rect 469864 6044 469916 6050
rect 469864 5986 469916 5992
rect 468484 5976 468536 5982
rect 468484 5918 468536 5924
rect 468668 3324 468720 3330
rect 468668 3266 468720 3272
rect 468680 480 468708 3266
rect 469876 480 469904 5986
rect 470612 490 470640 333610
rect 471992 16574 472020 336194
rect 475384 336184 475436 336190
rect 475384 336126 475436 336132
rect 486422 336152 486478 336161
rect 471992 16546 472296 16574
rect 470888 598 471100 626
rect 470888 490 470916 598
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 462 470916 490
rect 471072 480 471100 598
rect 472268 480 472296 16546
rect 473452 6112 473504 6118
rect 473452 6054 473504 6060
rect 473464 480 473492 6054
rect 474556 5976 474608 5982
rect 474556 5918 474608 5924
rect 474568 480 474596 5918
rect 475396 5574 475424 336126
rect 478880 336116 478932 336122
rect 486422 336087 486478 336096
rect 478880 336058 478932 336064
rect 477500 332172 477552 332178
rect 477500 332114 477552 332120
rect 477512 16574 477540 332114
rect 477512 16546 478184 16574
rect 476948 6792 477000 6798
rect 476948 6734 477000 6740
rect 475384 5568 475436 5574
rect 475384 5510 475436 5516
rect 475752 3392 475804 3398
rect 475752 3334 475804 3340
rect 475764 480 475792 3334
rect 476960 480 476988 6734
rect 478156 480 478184 16546
rect 478892 490 478920 336058
rect 483020 335300 483072 335306
rect 483020 335242 483072 335248
rect 481640 335232 481692 335238
rect 481640 335174 481692 335180
rect 481652 16574 481680 335174
rect 483032 16574 483060 335242
rect 485780 332104 485832 332110
rect 485780 332046 485832 332052
rect 485044 330880 485096 330886
rect 485044 330822 485096 330828
rect 481652 16546 482416 16574
rect 483032 16546 484072 16574
rect 481732 6724 481784 6730
rect 481732 6666 481784 6672
rect 480536 5568 480588 5574
rect 480536 5510 480588 5516
rect 479168 598 479380 626
rect 479168 490 479196 598
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 478892 462 479196 490
rect 479352 480 479380 598
rect 480548 480 480576 5510
rect 481744 480 481772 6666
rect 482388 490 482416 16546
rect 482664 598 482876 626
rect 482664 490 482692 598
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 462 482692 490
rect 482848 480 482876 598
rect 484044 480 484072 16546
rect 485056 3330 485084 330822
rect 485792 16574 485820 332046
rect 485792 16546 486372 16574
rect 485228 6656 485280 6662
rect 485228 6598 485280 6604
rect 485044 3324 485096 3330
rect 485044 3266 485096 3272
rect 485240 480 485268 6598
rect 486344 3482 486372 16546
rect 486436 5574 486464 336087
rect 497464 336048 497516 336054
rect 497464 335990 497516 335996
rect 504362 336016 504418 336025
rect 490012 335164 490064 335170
rect 490012 335106 490064 335112
rect 489184 332036 489236 332042
rect 489184 331978 489236 331984
rect 488816 6588 488868 6594
rect 488816 6530 488868 6536
rect 486424 5568 486476 5574
rect 486424 5510 486476 5516
rect 487620 5568 487672 5574
rect 487620 5510 487672 5516
rect 486344 3454 486464 3482
rect 486436 480 486464 3454
rect 487632 480 487660 5510
rect 488828 480 488856 6530
rect 489196 3398 489224 331978
rect 490024 16574 490052 335106
rect 492680 333600 492732 333606
rect 492680 333542 492732 333548
rect 492692 16574 492720 333542
rect 496820 331968 496872 331974
rect 496820 331910 496872 331916
rect 496832 16574 496860 331910
rect 490024 16546 490696 16574
rect 492692 16546 493088 16574
rect 496832 16546 497136 16574
rect 489184 3392 489236 3398
rect 489184 3334 489236 3340
rect 489920 3392 489972 3398
rect 489920 3334 489972 3340
rect 489932 480 489960 3334
rect 490668 490 490696 16546
rect 492312 6520 492364 6526
rect 492312 6462 492364 6468
rect 490944 598 491156 626
rect 490944 490 490972 598
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490668 462 490972 490
rect 491128 480 491156 598
rect 492324 480 492352 6462
rect 493060 490 493088 16546
rect 494704 8968 494756 8974
rect 494704 8910 494756 8916
rect 493336 598 493548 626
rect 493336 490 493364 598
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493060 462 493364 490
rect 493520 480 493548 598
rect 494716 480 494744 8910
rect 495900 6452 495952 6458
rect 495900 6394 495952 6400
rect 495912 480 495940 6394
rect 497108 480 497136 16546
rect 497476 5574 497504 335990
rect 504362 335951 504418 335960
rect 500960 335096 501012 335102
rect 500960 335038 501012 335044
rect 499580 330812 499632 330818
rect 499580 330754 499632 330760
rect 499592 16574 499620 330754
rect 500972 16574 501000 335038
rect 502984 333532 503036 333538
rect 502984 333474 503036 333480
rect 499592 16546 500632 16574
rect 500972 16546 501368 16574
rect 499396 6384 499448 6390
rect 499396 6326 499448 6332
rect 497464 5568 497516 5574
rect 497464 5510 497516 5516
rect 498200 5568 498252 5574
rect 498200 5510 498252 5516
rect 498212 480 498240 5510
rect 499408 480 499436 6326
rect 500604 480 500632 16546
rect 501340 490 501368 16546
rect 502892 6316 502944 6322
rect 502892 6258 502944 6264
rect 502904 3210 502932 6258
rect 502996 3330 503024 333474
rect 504376 5574 504404 335951
rect 507860 335028 507912 335034
rect 507860 334970 507912 334976
rect 506480 331900 506532 331906
rect 506480 331842 506532 331848
rect 506492 16574 506520 331842
rect 507872 16574 507900 334970
rect 512644 334960 512696 334966
rect 512644 334902 512696 334908
rect 510620 330744 510672 330750
rect 510620 330686 510672 330692
rect 510632 16574 510660 330686
rect 506492 16546 507256 16574
rect 507872 16546 508912 16574
rect 510632 16546 511304 16574
rect 506480 6248 506532 6254
rect 506480 6190 506532 6196
rect 504364 5568 504416 5574
rect 504364 5510 504416 5516
rect 505376 5568 505428 5574
rect 505376 5510 505428 5516
rect 502984 3324 503036 3330
rect 502984 3266 503036 3272
rect 504180 3324 504232 3330
rect 504180 3266 504232 3272
rect 502904 3182 503024 3210
rect 501616 598 501828 626
rect 501616 490 501644 598
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501340 462 501644 490
rect 501800 480 501828 598
rect 502996 480 503024 3182
rect 504192 480 504220 3266
rect 505388 480 505416 5510
rect 506492 480 506520 6190
rect 507228 490 507256 16546
rect 507504 598 507716 626
rect 507504 490 507532 598
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 462 507532 490
rect 507688 480 507716 598
rect 508884 480 508912 16546
rect 510068 6180 510120 6186
rect 510068 6122 510120 6128
rect 510080 480 510108 6122
rect 511276 480 511304 16546
rect 512460 4276 512512 4282
rect 512460 4218 512512 4224
rect 512472 480 512500 4218
rect 512656 3194 512684 334902
rect 520280 334892 520332 334898
rect 520280 334834 520332 334840
rect 515404 333464 515456 333470
rect 515404 333406 515456 333412
rect 514760 330676 514812 330682
rect 514760 330618 514812 330624
rect 512644 3188 512696 3194
rect 512644 3130 512696 3136
rect 513564 3188 513616 3194
rect 513564 3130 513616 3136
rect 513576 480 513604 3130
rect 514772 480 514800 330618
rect 515416 3330 515444 333406
rect 517520 330608 517572 330614
rect 517520 330550 517572 330556
rect 517532 16574 517560 330550
rect 519544 330540 519596 330546
rect 519544 330482 519596 330488
rect 519556 16574 519584 330482
rect 517532 16546 517928 16574
rect 519556 16546 519676 16574
rect 515956 4344 516008 4350
rect 515956 4286 516008 4292
rect 515404 3324 515456 3330
rect 515404 3266 515456 3272
rect 515968 480 515996 4286
rect 517152 3324 517204 3330
rect 517152 3266 517204 3272
rect 517164 480 517192 3266
rect 517900 490 517928 16546
rect 519544 4412 519596 4418
rect 519544 4354 519596 4360
rect 518176 598 518388 626
rect 518176 490 518204 598
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 462 518204 490
rect 518360 480 518388 598
rect 519556 480 519584 4354
rect 519648 3330 519676 16546
rect 519636 3324 519688 3330
rect 519636 3266 519688 3272
rect 520292 490 520320 334834
rect 526444 334824 526496 334830
rect 526444 334766 526496 334772
rect 522304 334756 522356 334762
rect 522304 334698 522356 334704
rect 522316 3330 522344 334698
rect 524420 329180 524472 329186
rect 524420 329122 524472 329128
rect 524432 16574 524460 329122
rect 524432 16546 525472 16574
rect 523040 4480 523092 4486
rect 523040 4422 523092 4428
rect 521844 3324 521896 3330
rect 521844 3266 521896 3272
rect 522304 3324 522356 3330
rect 522304 3266 522356 3272
rect 520568 598 520780 626
rect 520568 490 520596 598
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520292 462 520596 490
rect 520752 480 520780 598
rect 521856 480 521884 3266
rect 523052 480 523080 4422
rect 524236 3324 524288 3330
rect 524236 3266 524288 3272
rect 524248 480 524276 3266
rect 525444 480 525472 16546
rect 526456 3262 526484 334766
rect 528560 334688 528612 334694
rect 528560 334630 528612 334636
rect 526628 4548 526680 4554
rect 526628 4490 526680 4496
rect 526444 3256 526496 3262
rect 526444 3198 526496 3204
rect 526640 480 526668 4490
rect 527824 3256 527876 3262
rect 527824 3198 527876 3204
rect 527836 480 527864 3198
rect 528572 490 528600 334630
rect 540244 334620 540296 334626
rect 540244 334562 540296 334568
rect 530584 333396 530636 333402
rect 530584 333338 530636 333344
rect 530124 4616 530176 4622
rect 530124 4558 530176 4564
rect 528848 598 529060 626
rect 528848 490 528876 598
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528572 462 528876 490
rect 529032 480 529060 598
rect 530136 480 530164 4558
rect 530596 3398 530624 333338
rect 533344 333328 533396 333334
rect 533344 333270 533396 333276
rect 533356 3398 533384 333270
rect 538220 333260 538272 333266
rect 538220 333202 538272 333208
rect 535460 329112 535512 329118
rect 535460 329054 535512 329060
rect 535472 16574 535500 329054
rect 538232 16574 538260 333202
rect 535472 16546 536144 16574
rect 538232 16546 538444 16574
rect 533712 4684 533764 4690
rect 533712 4626 533764 4632
rect 530584 3392 530636 3398
rect 530584 3334 530636 3340
rect 531320 3392 531372 3398
rect 531320 3334 531372 3340
rect 533344 3392 533396 3398
rect 533344 3334 533396 3340
rect 531332 480 531360 3334
rect 532516 3324 532568 3330
rect 532516 3266 532568 3272
rect 532528 480 532556 3266
rect 533724 480 533752 4626
rect 534908 3392 534960 3398
rect 534908 3334 534960 3340
rect 534920 480 534948 3334
rect 536116 480 536144 16546
rect 537208 4752 537260 4758
rect 537208 4694 537260 4700
rect 537220 480 537248 4694
rect 538416 480 538444 16546
rect 540256 3398 540284 334562
rect 555436 313274 555464 459546
rect 556816 419490 556844 459614
rect 580264 458856 580316 458862
rect 580264 458798 580316 458804
rect 579802 458144 579858 458153
rect 579802 458079 579858 458088
rect 579816 456890 579844 458079
rect 579804 456884 579856 456890
rect 579804 456826 579856 456832
rect 580172 431928 580224 431934
rect 580172 431870 580224 431876
rect 580184 431633 580212 431870
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 556804 419484 556856 419490
rect 556804 419426 556856 419432
rect 580172 419484 580224 419490
rect 580172 419426 580224 419432
rect 580184 418305 580212 419426
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 579620 405680 579672 405686
rect 579620 405622 579672 405628
rect 579632 404977 579660 405622
rect 579618 404968 579674 404977
rect 579618 404903 579674 404912
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 579896 325644 579948 325650
rect 579896 325586 579948 325592
rect 579908 325281 579936 325586
rect 579894 325272 579950 325281
rect 579894 325207 579950 325216
rect 555424 313268 555476 313274
rect 555424 313210 555476 313216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580276 165889 580304 458798
rect 580262 165880 580318 165889
rect 580262 165815 580318 165824
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 545488 8220 545540 8226
rect 545488 8162 545540 8168
rect 540796 5500 540848 5506
rect 540796 5442 540848 5448
rect 539600 3392 539652 3398
rect 539600 3334 539652 3340
rect 540244 3392 540296 3398
rect 540244 3334 540296 3340
rect 539612 480 539640 3334
rect 540808 480 540836 5442
rect 544384 5432 544436 5438
rect 544384 5374 544436 5380
rect 543188 4072 543240 4078
rect 543188 4014 543240 4020
rect 541992 3392 542044 3398
rect 541992 3334 542044 3340
rect 542004 480 542032 3334
rect 543200 480 543228 4014
rect 544396 480 544424 5374
rect 545500 480 545528 8162
rect 549076 8152 549128 8158
rect 549076 8094 549128 8100
rect 547880 5364 547932 5370
rect 547880 5306 547932 5312
rect 546684 4004 546736 4010
rect 546684 3946 546736 3952
rect 546696 480 546724 3946
rect 547892 480 547920 5306
rect 549088 480 549116 8094
rect 552664 8084 552716 8090
rect 552664 8026 552716 8032
rect 551468 5296 551520 5302
rect 551468 5238 551520 5244
rect 550272 3936 550324 3942
rect 550272 3878 550324 3884
rect 550284 480 550312 3878
rect 551480 480 551508 5238
rect 552676 480 552704 8026
rect 556160 8016 556212 8022
rect 556160 7958 556212 7964
rect 554964 5228 555016 5234
rect 554964 5170 555016 5176
rect 553768 3868 553820 3874
rect 553768 3810 553820 3816
rect 553780 480 553808 3810
rect 554976 480 555004 5170
rect 556172 480 556200 7958
rect 559748 7948 559800 7954
rect 559748 7890 559800 7896
rect 558552 5160 558604 5166
rect 558552 5102 558604 5108
rect 557356 3800 557408 3806
rect 557356 3742 557408 3748
rect 557368 480 557396 3742
rect 558564 480 558592 5102
rect 559760 480 559788 7890
rect 563244 7880 563296 7886
rect 563244 7822 563296 7828
rect 562048 5092 562100 5098
rect 562048 5034 562100 5040
rect 560852 3732 560904 3738
rect 560852 3674 560904 3680
rect 560864 480 560892 3674
rect 562060 480 562088 5034
rect 563256 480 563284 7822
rect 566832 7812 566884 7818
rect 566832 7754 566884 7760
rect 565636 5024 565688 5030
rect 565636 4966 565688 4972
rect 564440 3664 564492 3670
rect 564440 3606 564492 3612
rect 564452 480 564480 3606
rect 565648 480 565676 4966
rect 566844 480 566872 7754
rect 570328 7744 570380 7750
rect 570328 7686 570380 7692
rect 569132 4956 569184 4962
rect 569132 4898 569184 4904
rect 568028 3596 568080 3602
rect 568028 3538 568080 3544
rect 568040 480 568068 3538
rect 569144 480 569172 4898
rect 570340 480 570368 7686
rect 573916 7676 573968 7682
rect 573916 7618 573968 7624
rect 572720 4888 572772 4894
rect 572720 4830 572772 4836
rect 571524 3528 571576 3534
rect 571524 3470 571576 3476
rect 571536 480 571564 3470
rect 572732 480 572760 4830
rect 573928 480 573956 7618
rect 577412 7608 577464 7614
rect 577412 7550 577464 7556
rect 576308 4820 576360 4826
rect 576308 4762 576360 4768
rect 575112 3460 575164 3466
rect 575112 3402 575164 3408
rect 575124 480 575152 3402
rect 576320 480 576348 4762
rect 577424 480 577452 7550
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 578606 3768 578662 3777
rect 578606 3703 578662 3712
rect 578620 480 578648 3703
rect 582194 3632 582250 3641
rect 582194 3567 582250 3576
rect 580998 3496 581054 3505
rect 580998 3431 581054 3440
rect 581012 480 581040 3431
rect 582208 480 582236 3567
rect 583390 3360 583446 3369
rect 583390 3295 583446 3304
rect 583404 480 583432 3295
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3146 658144 3202 658200
rect 2962 619112 3018 619168
rect 3330 606056 3386 606112
rect 3330 566888 3386 566944
rect 3330 553832 3386 553888
rect 3330 514820 3386 514856
rect 3330 514800 3332 514820
rect 3332 514800 3384 514820
rect 3384 514800 3386 514820
rect 3238 501744 3294 501800
rect 3514 671200 3570 671256
rect 3606 632032 3662 632088
rect 3698 579944 3754 580000
rect 3790 527856 3846 527912
rect 3974 475632 4030 475688
rect 3514 462576 3570 462632
rect 3330 449520 3386 449576
rect 3422 423544 3478 423600
rect 3422 410488 3478 410544
rect 3238 397432 3294 397488
rect 2778 371320 2834 371376
rect 3330 358400 3386 358456
rect 3146 345344 3202 345400
rect 43442 336368 43498 336424
rect 25502 336232 25558 336288
rect 18602 336096 18658 336152
rect 7562 335960 7618 336016
rect 3422 320048 3478 320104
rect 3422 319232 3478 319288
rect 3330 293800 3386 293856
rect 3330 293120 3386 293176
rect 3422 255176 3478 255232
rect 3422 254088 3478 254144
rect 3330 214920 3386 214976
rect 3422 202816 3478 202872
rect 3422 201864 3478 201920
rect 3422 164056 3478 164112
rect 3422 162832 3478 162888
rect 3422 137944 3478 138000
rect 3422 136720 3478 136776
rect 3422 111696 3478 111752
rect 3422 110608 3478 110664
rect 3422 85448 3478 85504
rect 3422 84632 3478 84688
rect 3330 59200 3386 59256
rect 3330 58520 3386 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3330 33088 3386 33144
rect 3330 32408 3386 32464
rect 3422 19352 3478 19408
rect 6458 3304 6514 3360
rect 15934 3576 15990 3632
rect 14738 3440 14794 3496
rect 24214 3712 24270 3768
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 237194 457272 237250 457328
rect 240782 457272 240838 457328
rect 242346 457272 242402 457328
rect 243910 457272 243966 457328
rect 245474 457272 245530 457328
rect 246946 457272 247002 457328
rect 248234 457272 248290 457328
rect 250258 457272 250314 457328
rect 251822 457272 251878 457328
rect 253386 457272 253442 457328
rect 256514 457272 256570 457328
rect 257526 457272 257582 457328
rect 259274 457272 259330 457328
rect 261298 457272 261354 457328
rect 262862 457272 262918 457328
rect 264518 457272 264574 457328
rect 266082 457272 266138 457328
rect 267554 457272 267610 457328
rect 269026 457272 269082 457328
rect 382278 457272 382334 457328
rect 384302 457272 384358 457328
rect 385406 457272 385462 457328
rect 387062 457272 387118 457328
rect 388626 457272 388682 457328
rect 390190 457272 390246 457328
rect 393502 457272 393558 457328
rect 394882 457272 394938 457328
rect 396538 457272 396594 457328
rect 398102 457272 398158 457328
rect 399666 457272 399722 457328
rect 401230 457272 401286 457328
rect 402978 457272 403034 457328
rect 404358 457272 404414 457328
rect 406014 457272 406070 457328
rect 409142 457272 409198 457328
rect 410706 457272 410762 457328
rect 412270 457272 412326 457328
rect 236274 335960 236330 336016
rect 238114 336096 238170 336152
rect 236274 3304 236330 3360
rect 241058 336368 241114 336424
rect 240690 336232 240746 336288
rect 238942 3576 238998 3632
rect 238850 3440 238906 3496
rect 241886 3712 241942 3768
rect 277122 3304 277178 3360
rect 283102 3440 283158 3496
rect 290186 3576 290242 3632
rect 294878 3712 294934 3768
rect 320270 3304 320326 3360
rect 321650 3440 321706 3496
rect 325974 3712 326030 3768
rect 324502 3576 324558 3632
rect 384670 336640 384726 336696
rect 385774 336096 385830 336152
rect 386878 336504 386934 336560
rect 387706 336232 387762 336288
rect 388994 336640 389050 336696
rect 391202 335960 391258 336016
rect 391938 336504 391994 336560
rect 417422 336232 417478 336288
rect 413926 3712 413982 3768
rect 415214 3576 415270 3632
rect 415122 3440 415178 3496
rect 415306 3304 415362 3360
rect 486422 336096 486478 336152
rect 504362 335960 504418 336016
rect 579802 458088 579858 458144
rect 580170 431568 580226 431624
rect 580170 418240 580226 418296
rect 579618 404912 579674 404968
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 580170 351872 580226 351928
rect 579894 325216 579950 325272
rect 580170 312024 580226 312080
rect 580262 165824 580318 165880
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
rect 578606 3712 578662 3768
rect 582194 3576 582250 3632
rect 580998 3440 581054 3496
rect 583390 3304 583446 3360
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3141 658202 3207 658205
rect -960 658200 3207 658202
rect -960 658144 3146 658200
rect 3202 658144 3207 658200
rect -960 658142 3207 658144
rect -960 658052 480 658142
rect 3141 658139 3207 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3601 632090 3667 632093
rect -960 632088 3667 632090
rect -960 632032 3606 632088
rect 3662 632032 3667 632088
rect -960 632030 3667 632032
rect -960 631940 480 632030
rect 3601 632027 3667 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 2957 619170 3023 619173
rect -960 619168 3023 619170
rect -960 619112 2962 619168
rect 3018 619112 3023 619168
rect -960 619110 3023 619112
rect -960 619020 480 619110
rect 2957 619107 3023 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3325 606114 3391 606117
rect -960 606112 3391 606114
rect -960 606056 3330 606112
rect 3386 606056 3391 606112
rect -960 606054 3391 606056
rect -960 605964 480 606054
rect 3325 606051 3391 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3693 580002 3759 580005
rect -960 580000 3759 580002
rect -960 579944 3698 580000
rect 3754 579944 3759 580000
rect -960 579942 3759 579944
rect -960 579852 480 579942
rect 3693 579939 3759 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3325 566946 3391 566949
rect -960 566944 3391 566946
rect -960 566888 3330 566944
rect 3386 566888 3391 566944
rect -960 566886 3391 566888
rect -960 566796 480 566886
rect 3325 566883 3391 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3785 527914 3851 527917
rect -960 527912 3851 527914
rect -960 527856 3790 527912
rect 3846 527856 3851 527912
rect -960 527854 3851 527856
rect -960 527764 480 527854
rect 3785 527851 3851 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3325 514858 3391 514861
rect -960 514856 3391 514858
rect -960 514800 3330 514856
rect 3386 514800 3391 514856
rect -960 514798 3391 514800
rect -960 514708 480 514798
rect 3325 514795 3391 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3233 501802 3299 501805
rect -960 501800 3299 501802
rect -960 501744 3238 501800
rect 3294 501744 3299 501800
rect -960 501742 3299 501744
rect -960 501652 480 501742
rect 3233 501739 3299 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3969 475690 4035 475693
rect -960 475688 4035 475690
rect -960 475632 3974 475688
rect 4030 475632 4035 475688
rect -960 475630 4035 475632
rect -960 475540 480 475630
rect 3969 475627 4035 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 579797 458146 579863 458149
rect 583520 458146 584960 458236
rect 579797 458144 584960 458146
rect 579797 458088 579802 458144
rect 579858 458088 584960 458144
rect 579797 458086 584960 458088
rect 579797 458083 579863 458086
rect 583520 457996 584960 458086
rect 237189 457332 237255 457333
rect 237189 457328 237236 457332
rect 237300 457330 237306 457332
rect 240777 457330 240843 457333
rect 241278 457330 241284 457332
rect 237189 457272 237194 457328
rect 237189 457268 237236 457272
rect 237300 457270 237346 457330
rect 240777 457328 241284 457330
rect 240777 457272 240782 457328
rect 240838 457272 241284 457328
rect 240777 457270 241284 457272
rect 237300 457268 237306 457270
rect 237189 457267 237255 457268
rect 240777 457267 240843 457270
rect 241278 457268 241284 457270
rect 241348 457268 241354 457332
rect 242341 457330 242407 457333
rect 242750 457330 242756 457332
rect 242341 457328 242756 457330
rect 242341 457272 242346 457328
rect 242402 457272 242756 457328
rect 242341 457270 242756 457272
rect 242341 457267 242407 457270
rect 242750 457268 242756 457270
rect 242820 457268 242826 457332
rect 243905 457330 243971 457333
rect 245469 457332 245535 457333
rect 244038 457330 244044 457332
rect 243905 457328 244044 457330
rect 243905 457272 243910 457328
rect 243966 457272 244044 457328
rect 243905 457270 244044 457272
rect 243905 457267 243971 457270
rect 244038 457268 244044 457270
rect 244108 457268 244114 457332
rect 245469 457328 245516 457332
rect 245580 457330 245586 457332
rect 245469 457272 245474 457328
rect 245469 457268 245516 457272
rect 245580 457270 245626 457330
rect 245580 457268 245586 457270
rect 246798 457268 246804 457332
rect 246868 457330 246874 457332
rect 246941 457330 247007 457333
rect 246868 457328 247007 457330
rect 246868 457272 246946 457328
rect 247002 457272 247007 457328
rect 246868 457270 247007 457272
rect 246868 457268 246874 457270
rect 245469 457267 245535 457268
rect 246941 457267 247007 457270
rect 248229 457332 248295 457333
rect 248229 457328 248276 457332
rect 248340 457330 248346 457332
rect 250253 457330 250319 457333
rect 251030 457330 251036 457332
rect 248229 457272 248234 457328
rect 248229 457268 248276 457272
rect 248340 457270 248386 457330
rect 250253 457328 251036 457330
rect 250253 457272 250258 457328
rect 250314 457272 251036 457328
rect 250253 457270 251036 457272
rect 248340 457268 248346 457270
rect 248229 457267 248295 457268
rect 250253 457267 250319 457270
rect 251030 457268 251036 457270
rect 251100 457268 251106 457332
rect 251817 457330 251883 457333
rect 252318 457330 252324 457332
rect 251817 457328 252324 457330
rect 251817 457272 251822 457328
rect 251878 457272 252324 457328
rect 251817 457270 252324 457272
rect 251817 457267 251883 457270
rect 252318 457268 252324 457270
rect 252388 457268 252394 457332
rect 253381 457330 253447 457333
rect 256509 457332 256575 457333
rect 253606 457330 253612 457332
rect 253381 457328 253612 457330
rect 253381 457272 253386 457328
rect 253442 457272 253612 457328
rect 253381 457270 253612 457272
rect 253381 457267 253447 457270
rect 253606 457268 253612 457270
rect 253676 457268 253682 457332
rect 256509 457328 256556 457332
rect 256620 457330 256626 457332
rect 256509 457272 256514 457328
rect 256509 457268 256556 457272
rect 256620 457270 256666 457330
rect 256620 457268 256626 457270
rect 257286 457268 257292 457332
rect 257356 457330 257362 457332
rect 257521 457330 257587 457333
rect 257356 457328 257587 457330
rect 257356 457272 257526 457328
rect 257582 457272 257587 457328
rect 257356 457270 257587 457272
rect 257356 457268 257362 457270
rect 256509 457267 256575 457268
rect 257521 457267 257587 457270
rect 259269 457332 259335 457333
rect 259269 457328 259316 457332
rect 259380 457330 259386 457332
rect 261293 457330 261359 457333
rect 262070 457330 262076 457332
rect 259269 457272 259274 457328
rect 259269 457268 259316 457272
rect 259380 457270 259426 457330
rect 261293 457328 262076 457330
rect 261293 457272 261298 457328
rect 261354 457272 262076 457328
rect 261293 457270 262076 457272
rect 259380 457268 259386 457270
rect 259269 457267 259335 457268
rect 261293 457267 261359 457270
rect 262070 457268 262076 457270
rect 262140 457268 262146 457332
rect 262857 457330 262923 457333
rect 263358 457330 263364 457332
rect 262857 457328 263364 457330
rect 262857 457272 262862 457328
rect 262918 457272 263364 457328
rect 262857 457270 263364 457272
rect 262857 457267 262923 457270
rect 263358 457268 263364 457270
rect 263428 457268 263434 457332
rect 264513 457330 264579 457333
rect 266077 457332 266143 457333
rect 267549 457332 267615 457333
rect 264646 457330 264652 457332
rect 264513 457328 264652 457330
rect 264513 457272 264518 457328
rect 264574 457272 264652 457328
rect 264513 457270 264652 457272
rect 264513 457267 264579 457270
rect 264646 457268 264652 457270
rect 264716 457268 264722 457332
rect 266077 457328 266124 457332
rect 266188 457330 266194 457332
rect 266077 457272 266082 457328
rect 266077 457268 266124 457272
rect 266188 457270 266234 457330
rect 267549 457328 267596 457332
rect 267660 457330 267666 457332
rect 267549 457272 267554 457328
rect 266188 457268 266194 457270
rect 267549 457268 267596 457272
rect 267660 457270 267706 457330
rect 267660 457268 267666 457270
rect 268878 457268 268884 457332
rect 268948 457330 268954 457332
rect 269021 457330 269087 457333
rect 382273 457332 382339 457333
rect 384297 457332 384363 457333
rect 382222 457330 382228 457332
rect 268948 457328 269087 457330
rect 268948 457272 269026 457328
rect 269082 457272 269087 457328
rect 268948 457270 269087 457272
rect 382182 457270 382228 457330
rect 382292 457328 382339 457332
rect 384246 457330 384252 457332
rect 382334 457272 382339 457328
rect 268948 457268 268954 457270
rect 266077 457267 266143 457268
rect 267549 457267 267615 457268
rect 269021 457267 269087 457270
rect 382222 457268 382228 457270
rect 382292 457268 382339 457272
rect 384206 457270 384252 457330
rect 384316 457328 384363 457332
rect 384358 457272 384363 457328
rect 384246 457268 384252 457270
rect 384316 457268 384363 457272
rect 384982 457268 384988 457332
rect 385052 457330 385058 457332
rect 385401 457330 385467 457333
rect 385052 457328 385467 457330
rect 385052 457272 385406 457328
rect 385462 457272 385467 457328
rect 385052 457270 385467 457272
rect 385052 457268 385058 457270
rect 382273 457267 382339 457268
rect 384297 457267 384363 457268
rect 385401 457267 385467 457270
rect 386454 457268 386460 457332
rect 386524 457330 386530 457332
rect 387057 457330 387123 457333
rect 386524 457328 387123 457330
rect 386524 457272 387062 457328
rect 387118 457272 387123 457328
rect 386524 457270 387123 457272
rect 386524 457268 386530 457270
rect 387057 457267 387123 457270
rect 387926 457268 387932 457332
rect 387996 457330 388002 457332
rect 388621 457330 388687 457333
rect 387996 457328 388687 457330
rect 387996 457272 388626 457328
rect 388682 457272 388687 457328
rect 387996 457270 388687 457272
rect 387996 457268 388002 457270
rect 388621 457267 388687 457270
rect 389214 457268 389220 457332
rect 389284 457330 389290 457332
rect 390185 457330 390251 457333
rect 393497 457332 393563 457333
rect 393446 457330 393452 457332
rect 389284 457328 390251 457330
rect 389284 457272 390190 457328
rect 390246 457272 390251 457328
rect 389284 457270 390251 457272
rect 393406 457270 393452 457330
rect 393516 457328 393563 457332
rect 393558 457272 393563 457328
rect 389284 457268 389290 457270
rect 390185 457267 390251 457270
rect 393446 457268 393452 457270
rect 393516 457268 393563 457272
rect 394734 457268 394740 457332
rect 394804 457330 394810 457332
rect 394877 457330 394943 457333
rect 394804 457328 394943 457330
rect 394804 457272 394882 457328
rect 394938 457272 394943 457328
rect 394804 457270 394943 457272
rect 394804 457268 394810 457270
rect 393497 457267 393563 457268
rect 394877 457267 394943 457270
rect 396206 457268 396212 457332
rect 396276 457330 396282 457332
rect 396533 457330 396599 457333
rect 396276 457328 396599 457330
rect 396276 457272 396538 457328
rect 396594 457272 396599 457328
rect 396276 457270 396599 457272
rect 396276 457268 396282 457270
rect 396533 457267 396599 457270
rect 397494 457268 397500 457332
rect 397564 457330 397570 457332
rect 398097 457330 398163 457333
rect 397564 457328 398163 457330
rect 397564 457272 398102 457328
rect 398158 457272 398163 457328
rect 397564 457270 398163 457272
rect 397564 457268 397570 457270
rect 398097 457267 398163 457270
rect 398782 457268 398788 457332
rect 398852 457330 398858 457332
rect 399661 457330 399727 457333
rect 398852 457328 399727 457330
rect 398852 457272 399666 457328
rect 399722 457272 399727 457328
rect 398852 457270 399727 457272
rect 398852 457268 398858 457270
rect 399661 457267 399727 457270
rect 400254 457268 400260 457332
rect 400324 457330 400330 457332
rect 401225 457330 401291 457333
rect 400324 457328 401291 457330
rect 400324 457272 401230 457328
rect 401286 457272 401291 457328
rect 400324 457270 401291 457272
rect 400324 457268 400330 457270
rect 401225 457267 401291 457270
rect 402973 457332 403039 457333
rect 404353 457332 404419 457333
rect 406009 457332 406075 457333
rect 402973 457328 403020 457332
rect 403084 457330 403090 457332
rect 404302 457330 404308 457332
rect 402973 457272 402978 457328
rect 402973 457268 403020 457272
rect 403084 457270 403130 457330
rect 404262 457270 404308 457330
rect 404372 457328 404419 457332
rect 405958 457330 405964 457332
rect 404414 457272 404419 457328
rect 403084 457268 403090 457270
rect 404302 457268 404308 457270
rect 404372 457268 404419 457272
rect 405918 457270 405964 457330
rect 406028 457328 406075 457332
rect 406070 457272 406075 457328
rect 405958 457268 405964 457270
rect 406028 457268 406075 457272
rect 408718 457268 408724 457332
rect 408788 457330 408794 457332
rect 409137 457330 409203 457333
rect 408788 457328 409203 457330
rect 408788 457272 409142 457328
rect 409198 457272 409203 457328
rect 408788 457270 409203 457272
rect 408788 457268 408794 457270
rect 402973 457267 403039 457268
rect 404353 457267 404419 457268
rect 406009 457267 406075 457268
rect 409137 457267 409203 457270
rect 409822 457268 409828 457332
rect 409892 457330 409898 457332
rect 410701 457330 410767 457333
rect 409892 457328 410767 457330
rect 409892 457272 410706 457328
rect 410762 457272 410767 457328
rect 409892 457270 410767 457272
rect 409892 457268 409898 457270
rect 410701 457267 410767 457270
rect 411294 457268 411300 457332
rect 411364 457330 411370 457332
rect 412265 457330 412331 457333
rect 411364 457328 412331 457330
rect 411364 457272 412270 457328
rect 412326 457272 412331 457328
rect 411364 457270 412331 457272
rect 411364 457268 411370 457270
rect 412265 457267 412331 457270
rect -960 449578 480 449668
rect 3325 449578 3391 449581
rect -960 449576 3391 449578
rect -960 449520 3330 449576
rect 3386 449520 3391 449576
rect -960 449518 3391 449520
rect -960 449428 480 449518
rect 3325 449515 3391 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3417 410546 3483 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect -960 410486 3483 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 579613 404970 579679 404973
rect 583520 404970 584960 405060
rect 579613 404968 584960 404970
rect 579613 404912 579618 404968
rect 579674 404912 584960 404968
rect 579613 404910 584960 404912
rect 579613 404907 579679 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3233 397490 3299 397493
rect -960 397488 3299 397490
rect -960 397432 3238 397488
rect 3294 397432 3299 397488
rect -960 397430 3299 397432
rect -960 397340 480 397430
rect 3233 397427 3299 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 2773 371378 2839 371381
rect -960 371376 2839 371378
rect -960 371320 2778 371376
rect 2834 371320 2839 371376
rect -960 371318 2839 371320
rect -960 371228 480 371318
rect 2773 371315 2839 371318
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3141 345402 3207 345405
rect -960 345400 3207 345402
rect -960 345344 3146 345400
rect 3202 345344 3207 345400
rect -960 345342 3207 345344
rect -960 345252 480 345342
rect 3141 345339 3207 345342
rect 583520 338452 584960 338692
rect 384665 336698 384731 336701
rect 388989 336698 389055 336701
rect 384665 336696 389055 336698
rect 384665 336640 384670 336696
rect 384726 336640 388994 336696
rect 389050 336640 389055 336696
rect 384665 336638 389055 336640
rect 384665 336635 384731 336638
rect 388989 336635 389055 336638
rect 386873 336562 386939 336565
rect 391933 336562 391999 336565
rect 386873 336560 391999 336562
rect 386873 336504 386878 336560
rect 386934 336504 391938 336560
rect 391994 336504 391999 336560
rect 386873 336502 391999 336504
rect 386873 336499 386939 336502
rect 391933 336499 391999 336502
rect 43437 336426 43503 336429
rect 241053 336426 241119 336429
rect 43437 336424 241119 336426
rect 43437 336368 43442 336424
rect 43498 336368 241058 336424
rect 241114 336368 241119 336424
rect 43437 336366 241119 336368
rect 43437 336363 43503 336366
rect 241053 336363 241119 336366
rect 25497 336290 25563 336293
rect 240685 336290 240751 336293
rect 25497 336288 240751 336290
rect 25497 336232 25502 336288
rect 25558 336232 240690 336288
rect 240746 336232 240751 336288
rect 25497 336230 240751 336232
rect 25497 336227 25563 336230
rect 240685 336227 240751 336230
rect 387701 336290 387767 336293
rect 417417 336290 417483 336293
rect 387701 336288 417483 336290
rect 387701 336232 387706 336288
rect 387762 336232 417422 336288
rect 417478 336232 417483 336288
rect 387701 336230 417483 336232
rect 387701 336227 387767 336230
rect 417417 336227 417483 336230
rect 18597 336154 18663 336157
rect 238109 336154 238175 336157
rect 18597 336152 238175 336154
rect 18597 336096 18602 336152
rect 18658 336096 238114 336152
rect 238170 336096 238175 336152
rect 18597 336094 238175 336096
rect 18597 336091 18663 336094
rect 238109 336091 238175 336094
rect 385769 336154 385835 336157
rect 486417 336154 486483 336157
rect 385769 336152 486483 336154
rect 385769 336096 385774 336152
rect 385830 336096 486422 336152
rect 486478 336096 486483 336152
rect 385769 336094 486483 336096
rect 385769 336091 385835 336094
rect 486417 336091 486483 336094
rect 7557 336018 7623 336021
rect 236269 336018 236335 336021
rect 7557 336016 236335 336018
rect 7557 335960 7562 336016
rect 7618 335960 236274 336016
rect 236330 335960 236335 336016
rect 7557 335958 236335 335960
rect 7557 335955 7623 335958
rect 236269 335955 236335 335958
rect 391197 336018 391263 336021
rect 504357 336018 504423 336021
rect 391197 336016 504423 336018
rect 391197 335960 391202 336016
rect 391258 335960 504362 336016
rect 504418 335960 504423 336016
rect 391197 335958 504423 335960
rect 391197 335955 391263 335958
rect 504357 335955 504423 335958
rect -960 332196 480 332436
rect 579889 325274 579955 325277
rect 583520 325274 584960 325364
rect 579889 325272 584960 325274
rect 579889 325216 579894 325272
rect 579950 325216 584960 325272
rect 579889 325214 584960 325216
rect 579889 325211 579955 325214
rect 583520 325124 584960 325214
rect 3417 320106 3483 320109
rect 382222 320106 382228 320108
rect 3417 320104 382228 320106
rect 3417 320048 3422 320104
rect 3478 320048 382228 320104
rect 3417 320046 382228 320048
rect 3417 320043 3483 320046
rect 382222 320044 382228 320046
rect 382292 320044 382298 320108
rect -960 319290 480 319380
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect 384982 306370 384988 306372
rect -960 306234 480 306324
rect 6870 306310 384988 306370
rect 6870 306234 6930 306310
rect 384982 306308 384988 306310
rect 385052 306308 385058 306372
rect -960 306174 6930 306234
rect -960 306084 480 306174
rect 583520 298754 584960 298844
rect 583342 298694 584960 298754
rect 583342 298618 583402 298694
rect 583520 298618 584960 298694
rect 583342 298604 584960 298618
rect 583342 298558 583586 298604
rect 268878 298148 268884 298212
rect 268948 298210 268954 298212
rect 583526 298210 583586 298558
rect 268948 298150 583586 298210
rect 268948 298148 268954 298150
rect 3325 293858 3391 293861
rect 384246 293858 384252 293860
rect 3325 293856 384252 293858
rect 3325 293800 3330 293856
rect 3386 293800 384252 293856
rect 3325 293798 384252 293800
rect 3325 293795 3391 293798
rect 384246 293796 384252 293798
rect 384316 293796 384322 293860
rect -960 293178 480 293268
rect 3325 293178 3391 293181
rect -960 293176 3391 293178
rect -960 293120 3330 293176
rect 3386 293120 3391 293176
rect -960 293118 3391 293120
rect -960 293028 480 293118
rect 3325 293115 3391 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272234 584960 272324
rect 567150 272174 584960 272234
rect 266118 271900 266124 271964
rect 266188 271962 266194 271964
rect 567150 271962 567210 272174
rect 583520 272084 584960 272174
rect 266188 271902 567210 271962
rect 266188 271900 266194 271902
rect 386454 267746 386460 267748
rect 430 267686 386460 267746
rect 430 267474 490 267686
rect 386454 267684 386460 267686
rect 386524 267684 386530 267748
rect 430 267414 674 267474
rect -960 267202 480 267292
rect 614 267202 674 267414
rect -960 267142 674 267202
rect -960 267052 480 267142
rect 583520 258906 584960 258996
rect 583342 258846 584960 258906
rect 583342 258770 583402 258846
rect 583520 258770 584960 258846
rect 583342 258756 584960 258770
rect 583342 258710 583586 258756
rect 267590 258028 267596 258092
rect 267660 258090 267666 258092
rect 267660 258030 267842 258090
rect 267660 258028 267666 258030
rect 267782 257954 267842 258030
rect 583526 257954 583586 258710
rect 267782 257894 583586 257954
rect 3417 255234 3483 255237
rect 389214 255234 389220 255236
rect 3417 255232 389220 255234
rect 3417 255176 3422 255232
rect 3478 255176 389220 255232
rect 3417 255174 389220 255176
rect 3417 255171 3483 255174
rect 389214 255172 389220 255174
rect 389284 255172 389290 255236
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 583520 245578 584960 245668
rect 583342 245518 584960 245578
rect 583342 245442 583402 245518
rect 583520 245442 584960 245518
rect 583342 245428 584960 245442
rect 583342 245382 583586 245428
rect 264646 244292 264652 244356
rect 264716 244354 264722 244356
rect 583526 244354 583586 245382
rect 264716 244294 583586 244354
rect 264716 244292 264722 244294
rect 388110 241498 388116 241500
rect 6870 241438 388116 241498
rect -960 241090 480 241180
rect 6870 241090 6930 241438
rect 388110 241436 388116 241438
rect 388180 241436 388186 241500
rect -960 241030 6930 241090
rect -960 240940 480 241030
rect 583520 232386 584960 232476
rect 583342 232326 584960 232386
rect 583342 232250 583402 232326
rect 583520 232250 584960 232326
rect 583342 232236 584960 232250
rect 583342 232190 583586 232236
rect 262070 231916 262076 231980
rect 262140 231978 262146 231980
rect 583526 231978 583586 232190
rect 262140 231918 583586 231978
rect 262140 231916 262146 231918
rect -960 227884 480 228124
rect 583520 219058 584960 219148
rect 583342 218998 584960 219058
rect 583342 218922 583402 218998
rect 583520 218922 584960 218998
rect 583342 218908 584960 218922
rect 583342 218862 583586 218908
rect 263358 218044 263364 218108
rect 263428 218106 263434 218108
rect 583526 218106 583586 218862
rect 263428 218046 583586 218106
rect 263428 218044 263434 218046
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 259310 205668 259316 205732
rect 259380 205730 259386 205732
rect 583520 205730 584960 205820
rect 259380 205670 584960 205730
rect 259380 205668 259386 205670
rect 583520 205580 584960 205670
rect 3417 202874 3483 202877
rect 394734 202874 394740 202876
rect 3417 202872 394740 202874
rect 3417 202816 3422 202872
rect 3478 202816 394740 202872
rect 3417 202814 394740 202816
rect 3417 202811 3483 202814
rect 394734 202812 394740 202814
rect 394804 202812 394810 202876
rect -960 201922 480 202012
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 583520 192538 584960 192628
rect 583342 192478 584960 192538
rect 583342 192402 583402 192478
rect 583520 192402 584960 192478
rect 583342 192388 584960 192402
rect 583342 192342 583586 192388
rect 256550 191796 256556 191860
rect 256620 191858 256626 191860
rect 583526 191858 583586 192342
rect 256620 191798 583586 191858
rect 256620 191796 256626 191798
rect 393078 189002 393084 189004
rect -960 188866 480 188956
rect 6870 188942 393084 189002
rect 6870 188866 6930 188942
rect 393078 188940 393084 188942
rect 393148 188940 393154 189004
rect -960 188806 6930 188866
rect -960 188716 480 188806
rect 583520 179210 584960 179300
rect 583342 179150 584960 179210
rect 583342 179074 583402 179150
rect 583520 179074 584960 179150
rect 583342 179060 584960 179074
rect 583342 179014 583586 179060
rect 257286 178060 257292 178124
rect 257356 178122 257362 178124
rect 583526 178122 583586 179014
rect 257356 178062 583586 178122
rect 257356 178060 257362 178062
rect -960 175796 480 176036
rect 580257 165882 580323 165885
rect 583520 165882 584960 165972
rect 580257 165880 584960 165882
rect 580257 165824 580262 165880
rect 580318 165824 584960 165880
rect 580257 165822 584960 165824
rect 580257 165819 580323 165822
rect 583520 165732 584960 165822
rect 3417 164114 3483 164117
rect 396206 164114 396212 164116
rect 3417 164112 396212 164114
rect 3417 164056 3422 164112
rect 3478 164056 396212 164112
rect 3417 164054 396212 164056
rect 3417 164051 3483 164054
rect 396206 164052 396212 164054
rect 396276 164052 396282 164116
rect -960 162890 480 162980
rect 3417 162890 3483 162893
rect -960 162888 3483 162890
rect -960 162832 3422 162888
rect 3478 162832 3483 162888
rect -960 162830 3483 162832
rect -960 162740 480 162830
rect 3417 162827 3483 162830
rect 583520 152690 584960 152780
rect 583342 152630 584960 152690
rect 583342 152554 583402 152630
rect 583520 152554 584960 152630
rect 583342 152540 584960 152554
rect 583342 152494 583586 152540
rect 252318 151812 252324 151876
rect 252388 151874 252394 151876
rect 583526 151874 583586 152494
rect 252388 151814 583586 151874
rect 252388 151812 252394 151814
rect 398782 150378 398788 150380
rect 430 150318 398788 150378
rect 430 150106 490 150318
rect 398782 150316 398788 150318
rect 398852 150316 398858 150380
rect 430 150046 674 150106
rect -960 149834 480 149924
rect 614 149834 674 150046
rect -960 149774 674 149834
rect -960 149684 480 149774
rect 583520 139362 584960 139452
rect 583342 139302 584960 139362
rect 583342 139226 583402 139302
rect 583520 139226 584960 139302
rect 583342 139212 584960 139226
rect 583342 139166 583586 139212
rect 253606 138076 253612 138140
rect 253676 138138 253682 138140
rect 583526 138138 583586 139166
rect 253676 138078 583586 138138
rect 253676 138076 253682 138078
rect 3417 138002 3483 138005
rect 397494 138002 397500 138004
rect 3417 138000 397500 138002
rect 3417 137944 3422 138000
rect 3478 137944 397500 138000
rect 3417 137942 397500 137944
rect 3417 137939 3483 137942
rect 397494 137940 397500 137942
rect 397564 137940 397570 138004
rect -960 136778 480 136868
rect 3417 136778 3483 136781
rect -960 136776 3483 136778
rect -960 136720 3422 136776
rect 3478 136720 3483 136776
rect -960 136718 3483 136720
rect -960 136628 480 136718
rect 3417 136715 3483 136718
rect 583520 126034 584960 126124
rect 583342 125974 584960 126034
rect 583342 125898 583402 125974
rect 583520 125898 584960 125974
rect 583342 125884 584960 125898
rect 583342 125838 583586 125884
rect 251030 125564 251036 125628
rect 251100 125626 251106 125628
rect 583526 125626 583586 125838
rect 251100 125566 583586 125626
rect 251100 125564 251106 125566
rect -960 123572 480 123812
rect 583520 112842 584960 112932
rect 583342 112782 584960 112842
rect 583342 112706 583402 112782
rect 583520 112706 584960 112782
rect 583342 112692 584960 112706
rect 583342 112646 583586 112692
rect 246798 111828 246804 111892
rect 246868 111890 246874 111892
rect 583526 111890 583586 112646
rect 246868 111830 583586 111890
rect 246868 111828 246874 111830
rect 3417 111754 3483 111757
rect 400254 111754 400260 111756
rect 3417 111752 400260 111754
rect 3417 111696 3422 111752
rect 3478 111696 400260 111752
rect 3417 111694 400260 111696
rect 3417 111691 3483 111694
rect 400254 111692 400260 111694
rect 400324 111692 400330 111756
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 248270 99452 248276 99516
rect 248340 99514 248346 99516
rect 583520 99514 584960 99604
rect 248340 99454 584960 99514
rect 248340 99452 248346 99454
rect 583520 99364 584960 99454
rect 404302 97882 404308 97884
rect 6870 97822 404308 97882
rect -960 97610 480 97700
rect 6870 97610 6930 97822
rect 404302 97820 404308 97822
rect 404372 97820 404378 97884
rect -960 97550 6930 97610
rect -960 97460 480 97550
rect 583520 86186 584960 86276
rect 583342 86126 584960 86186
rect 583342 86050 583402 86126
rect 583520 86050 584960 86126
rect 583342 86036 584960 86050
rect 583342 85990 583586 86036
rect 245510 85580 245516 85644
rect 245580 85642 245586 85644
rect 583526 85642 583586 85990
rect 245580 85582 583586 85642
rect 245580 85580 245586 85582
rect 3417 85506 3483 85509
rect 403014 85506 403020 85508
rect 3417 85504 403020 85506
rect 3417 85448 3422 85504
rect 3478 85448 403020 85504
rect 3417 85446 403020 85448
rect 3417 85443 3483 85446
rect 403014 85444 403020 85446
rect 403084 85444 403090 85508
rect -960 84690 480 84780
rect 3417 84690 3483 84693
rect -960 84688 3483 84690
rect -960 84632 3422 84688
rect 3478 84632 3483 84688
rect -960 84630 3483 84632
rect -960 84540 480 84630
rect 3417 84627 3483 84630
rect 583520 72994 584960 73084
rect 583342 72934 584960 72994
rect 583342 72858 583402 72934
rect 583520 72858 584960 72934
rect 583342 72844 584960 72858
rect 583342 72798 583586 72844
rect 242750 71844 242756 71908
rect 242820 71906 242826 71908
rect 583526 71906 583586 72798
rect 242820 71846 583586 71906
rect 242820 71844 242826 71846
rect 405958 71770 405964 71772
rect -960 71634 480 71724
rect 6870 71710 405964 71770
rect 6870 71634 6930 71710
rect 405958 71708 405964 71710
rect 406028 71708 406034 71772
rect -960 71574 6930 71634
rect -960 71484 480 71574
rect 583520 59666 584960 59756
rect 567150 59606 584960 59666
rect 244038 59332 244044 59396
rect 244108 59394 244114 59396
rect 567150 59394 567210 59606
rect 583520 59516 584960 59606
rect 244108 59334 567210 59394
rect 244108 59332 244114 59334
rect 3325 59258 3391 59261
rect 408718 59258 408724 59260
rect 3325 59256 408724 59258
rect 3325 59200 3330 59256
rect 3386 59200 408724 59256
rect 3325 59198 408724 59200
rect 3325 59195 3391 59198
rect 408718 59196 408724 59198
rect 408788 59196 408794 59260
rect -960 58578 480 58668
rect 3325 58578 3391 58581
rect -960 58576 3391 58578
rect -960 58520 3330 58576
rect 3386 58520 3391 58576
rect -960 58518 3391 58520
rect -960 58428 480 58518
rect 3325 58515 3391 58518
rect 583520 46338 584960 46428
rect 583342 46278 584960 46338
rect 583342 46202 583402 46278
rect 583520 46202 584960 46278
rect 583342 46188 584960 46202
rect 583342 46142 583586 46188
rect -960 45522 480 45612
rect 241278 45596 241284 45660
rect 241348 45658 241354 45660
rect 583526 45658 583586 46142
rect 241348 45598 583586 45658
rect 241348 45596 241354 45598
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 3325 33146 3391 33149
rect 409822 33146 409828 33148
rect 3325 33144 409828 33146
rect 3325 33088 3330 33144
rect 3386 33088 409828 33144
rect 3325 33086 409828 33088
rect 3325 33083 3391 33086
rect 409822 33084 409828 33086
rect 409892 33084 409898 33148
rect 583520 33146 584960 33236
rect 583342 33086 584960 33146
rect 583342 33010 583402 33086
rect 583520 33010 584960 33086
rect 583342 32996 584960 33010
rect 583342 32950 583586 32996
rect -960 32466 480 32556
rect 3325 32466 3391 32469
rect -960 32464 3391 32466
rect -960 32408 3330 32464
rect 3386 32408 3391 32464
rect -960 32406 3391 32408
rect -960 32316 480 32406
rect 3325 32403 3391 32406
rect 237230 31724 237236 31788
rect 237300 31786 237306 31788
rect 583526 31786 583586 32950
rect 237300 31726 583586 31786
rect 237300 31724 237306 31726
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 411294 6898 411300 6900
rect 6870 6838 411300 6898
rect -960 6490 480 6580
rect 6870 6490 6930 6838
rect 411294 6836 411300 6838
rect 411364 6836 411370 6900
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect -960 6430 6930 6490
rect 583520 6476 584960 6566
rect -960 6340 480 6430
rect 24209 3770 24275 3773
rect 241881 3770 241947 3773
rect 24209 3768 241947 3770
rect 24209 3712 24214 3768
rect 24270 3712 241886 3768
rect 241942 3712 241947 3768
rect 24209 3710 241947 3712
rect 24209 3707 24275 3710
rect 241881 3707 241947 3710
rect 294873 3770 294939 3773
rect 325969 3770 326035 3773
rect 294873 3768 326035 3770
rect 294873 3712 294878 3768
rect 294934 3712 325974 3768
rect 326030 3712 326035 3768
rect 294873 3710 326035 3712
rect 294873 3707 294939 3710
rect 325969 3707 326035 3710
rect 413921 3770 413987 3773
rect 578601 3770 578667 3773
rect 413921 3768 578667 3770
rect 413921 3712 413926 3768
rect 413982 3712 578606 3768
rect 578662 3712 578667 3768
rect 413921 3710 578667 3712
rect 413921 3707 413987 3710
rect 578601 3707 578667 3710
rect 15929 3634 15995 3637
rect 238937 3634 239003 3637
rect 15929 3632 239003 3634
rect 15929 3576 15934 3632
rect 15990 3576 238942 3632
rect 238998 3576 239003 3632
rect 15929 3574 239003 3576
rect 15929 3571 15995 3574
rect 238937 3571 239003 3574
rect 290181 3634 290247 3637
rect 324497 3634 324563 3637
rect 290181 3632 324563 3634
rect 290181 3576 290186 3632
rect 290242 3576 324502 3632
rect 324558 3576 324563 3632
rect 290181 3574 324563 3576
rect 290181 3571 290247 3574
rect 324497 3571 324563 3574
rect 415209 3634 415275 3637
rect 582189 3634 582255 3637
rect 415209 3632 582255 3634
rect 415209 3576 415214 3632
rect 415270 3576 582194 3632
rect 582250 3576 582255 3632
rect 415209 3574 582255 3576
rect 415209 3571 415275 3574
rect 582189 3571 582255 3574
rect 14733 3498 14799 3501
rect 238845 3498 238911 3501
rect 14733 3496 238911 3498
rect 14733 3440 14738 3496
rect 14794 3440 238850 3496
rect 238906 3440 238911 3496
rect 14733 3438 238911 3440
rect 14733 3435 14799 3438
rect 238845 3435 238911 3438
rect 283097 3498 283163 3501
rect 321645 3498 321711 3501
rect 283097 3496 321711 3498
rect 283097 3440 283102 3496
rect 283158 3440 321650 3496
rect 321706 3440 321711 3496
rect 283097 3438 321711 3440
rect 283097 3435 283163 3438
rect 321645 3435 321711 3438
rect 415117 3498 415183 3501
rect 580993 3498 581059 3501
rect 415117 3496 581059 3498
rect 415117 3440 415122 3496
rect 415178 3440 580998 3496
rect 581054 3440 581059 3496
rect 415117 3438 581059 3440
rect 415117 3435 415183 3438
rect 580993 3435 581059 3438
rect 6453 3362 6519 3365
rect 236269 3362 236335 3365
rect 6453 3360 236335 3362
rect 6453 3304 6458 3360
rect 6514 3304 236274 3360
rect 236330 3304 236335 3360
rect 6453 3302 236335 3304
rect 6453 3299 6519 3302
rect 236269 3299 236335 3302
rect 277117 3362 277183 3365
rect 320265 3362 320331 3365
rect 277117 3360 320331 3362
rect 277117 3304 277122 3360
rect 277178 3304 320270 3360
rect 320326 3304 320331 3360
rect 277117 3302 320331 3304
rect 277117 3299 277183 3302
rect 320265 3299 320331 3302
rect 415301 3362 415367 3365
rect 583385 3362 583451 3365
rect 415301 3360 583451 3362
rect 415301 3304 415306 3360
rect 415362 3304 583390 3360
rect 583446 3304 583451 3360
rect 415301 3302 583451 3304
rect 415301 3299 415367 3302
rect 583385 3299 583451 3302
<< via3 >>
rect 237236 457328 237300 457332
rect 237236 457272 237250 457328
rect 237250 457272 237300 457328
rect 237236 457268 237300 457272
rect 241284 457268 241348 457332
rect 242756 457268 242820 457332
rect 244044 457268 244108 457332
rect 245516 457328 245580 457332
rect 245516 457272 245530 457328
rect 245530 457272 245580 457328
rect 245516 457268 245580 457272
rect 246804 457268 246868 457332
rect 248276 457328 248340 457332
rect 248276 457272 248290 457328
rect 248290 457272 248340 457328
rect 248276 457268 248340 457272
rect 251036 457268 251100 457332
rect 252324 457268 252388 457332
rect 253612 457268 253676 457332
rect 256556 457328 256620 457332
rect 256556 457272 256570 457328
rect 256570 457272 256620 457328
rect 256556 457268 256620 457272
rect 257292 457268 257356 457332
rect 259316 457328 259380 457332
rect 259316 457272 259330 457328
rect 259330 457272 259380 457328
rect 259316 457268 259380 457272
rect 262076 457268 262140 457332
rect 263364 457268 263428 457332
rect 264652 457268 264716 457332
rect 266124 457328 266188 457332
rect 266124 457272 266138 457328
rect 266138 457272 266188 457328
rect 266124 457268 266188 457272
rect 267596 457328 267660 457332
rect 267596 457272 267610 457328
rect 267610 457272 267660 457328
rect 267596 457268 267660 457272
rect 268884 457268 268948 457332
rect 382228 457328 382292 457332
rect 382228 457272 382278 457328
rect 382278 457272 382292 457328
rect 382228 457268 382292 457272
rect 384252 457328 384316 457332
rect 384252 457272 384302 457328
rect 384302 457272 384316 457328
rect 384252 457268 384316 457272
rect 384988 457268 385052 457332
rect 386460 457268 386524 457332
rect 387932 457268 387996 457332
rect 389220 457268 389284 457332
rect 393452 457328 393516 457332
rect 393452 457272 393502 457328
rect 393502 457272 393516 457328
rect 393452 457268 393516 457272
rect 394740 457268 394804 457332
rect 396212 457268 396276 457332
rect 397500 457268 397564 457332
rect 398788 457268 398852 457332
rect 400260 457268 400324 457332
rect 403020 457328 403084 457332
rect 403020 457272 403034 457328
rect 403034 457272 403084 457328
rect 403020 457268 403084 457272
rect 404308 457328 404372 457332
rect 404308 457272 404358 457328
rect 404358 457272 404372 457328
rect 404308 457268 404372 457272
rect 405964 457328 406028 457332
rect 405964 457272 406014 457328
rect 406014 457272 406028 457328
rect 405964 457268 406028 457272
rect 408724 457268 408788 457332
rect 409828 457268 409892 457332
rect 411300 457268 411364 457332
rect 382228 320044 382292 320108
rect 384988 306308 385052 306372
rect 268884 298148 268948 298212
rect 384252 293796 384316 293860
rect 266124 271900 266188 271964
rect 386460 267684 386524 267748
rect 267596 258028 267660 258092
rect 389220 255172 389284 255236
rect 264652 244292 264716 244356
rect 388116 241436 388180 241500
rect 262076 231916 262140 231980
rect 263364 218044 263428 218108
rect 259316 205668 259380 205732
rect 394740 202812 394804 202876
rect 256556 191796 256620 191860
rect 393084 188940 393148 189004
rect 257292 178060 257356 178124
rect 396212 164052 396276 164116
rect 252324 151812 252388 151876
rect 398788 150316 398852 150380
rect 253612 138076 253676 138140
rect 397500 137940 397564 138004
rect 251036 125564 251100 125628
rect 246804 111828 246868 111892
rect 400260 111692 400324 111756
rect 248276 99452 248340 99516
rect 404308 97820 404372 97884
rect 245516 85580 245580 85644
rect 403020 85444 403084 85508
rect 242756 71844 242820 71908
rect 405964 71708 406028 71772
rect 244044 59332 244108 59396
rect 408724 59196 408788 59260
rect 241284 45596 241348 45660
rect 409828 33084 409892 33148
rect 237236 31724 237300 31788
rect 411300 6836 411364 6900
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711002 -8694 711558
rect -8138 711002 -8106 711558
rect -8726 680614 -8106 711002
rect -8726 680058 -8694 680614
rect -8138 680058 -8106 680614
rect -8726 644614 -8106 680058
rect -8726 644058 -8694 644614
rect -8138 644058 -8106 644614
rect -8726 608614 -8106 644058
rect -8726 608058 -8694 608614
rect -8138 608058 -8106 608614
rect -8726 572614 -8106 608058
rect -8726 572058 -8694 572614
rect -8138 572058 -8106 572614
rect -8726 536614 -8106 572058
rect -8726 536058 -8694 536614
rect -8138 536058 -8106 536614
rect -8726 500614 -8106 536058
rect -8726 500058 -8694 500614
rect -8138 500058 -8106 500614
rect -8726 464614 -8106 500058
rect -8726 464058 -8694 464614
rect -8138 464058 -8106 464614
rect -8726 428614 -8106 464058
rect -8726 428058 -8694 428614
rect -8138 428058 -8106 428614
rect -8726 392614 -8106 428058
rect -8726 392058 -8694 392614
rect -8138 392058 -8106 392614
rect -8726 356614 -8106 392058
rect -8726 356058 -8694 356614
rect -8138 356058 -8106 356614
rect -8726 320614 -8106 356058
rect -8726 320058 -8694 320614
rect -8138 320058 -8106 320614
rect -8726 284614 -8106 320058
rect -8726 284058 -8694 284614
rect -8138 284058 -8106 284614
rect -8726 248614 -8106 284058
rect -8726 248058 -8694 248614
rect -8138 248058 -8106 248614
rect -8726 212614 -8106 248058
rect -8726 212058 -8694 212614
rect -8138 212058 -8106 212614
rect -8726 176614 -8106 212058
rect -8726 176058 -8694 176614
rect -8138 176058 -8106 176614
rect -8726 140614 -8106 176058
rect -8726 140058 -8694 140614
rect -8138 140058 -8106 140614
rect -8726 104614 -8106 140058
rect -8726 104058 -8694 104614
rect -8138 104058 -8106 104614
rect -8726 68614 -8106 104058
rect -8726 68058 -8694 68614
rect -8138 68058 -8106 68614
rect -8726 32614 -8106 68058
rect -8726 32058 -8694 32614
rect -8138 32058 -8106 32614
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710042 -7734 710598
rect -7178 710042 -7146 710598
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710042 12986 710598
rect 13542 710042 13574 710598
rect -7766 698058 -7734 698614
rect -7178 698058 -7146 698614
rect -7766 662614 -7146 698058
rect -7766 662058 -7734 662614
rect -7178 662058 -7146 662614
rect -7766 626614 -7146 662058
rect -7766 626058 -7734 626614
rect -7178 626058 -7146 626614
rect -7766 590614 -7146 626058
rect -7766 590058 -7734 590614
rect -7178 590058 -7146 590614
rect -7766 554614 -7146 590058
rect -7766 554058 -7734 554614
rect -7178 554058 -7146 554614
rect -7766 518614 -7146 554058
rect -7766 518058 -7734 518614
rect -7178 518058 -7146 518614
rect -7766 482614 -7146 518058
rect -7766 482058 -7734 482614
rect -7178 482058 -7146 482614
rect -7766 446614 -7146 482058
rect -7766 446058 -7734 446614
rect -7178 446058 -7146 446614
rect -7766 410614 -7146 446058
rect -7766 410058 -7734 410614
rect -7178 410058 -7146 410614
rect -7766 374614 -7146 410058
rect -7766 374058 -7734 374614
rect -7178 374058 -7146 374614
rect -7766 338614 -7146 374058
rect -7766 338058 -7734 338614
rect -7178 338058 -7146 338614
rect -7766 302614 -7146 338058
rect -7766 302058 -7734 302614
rect -7178 302058 -7146 302614
rect -7766 266614 -7146 302058
rect -7766 266058 -7734 266614
rect -7178 266058 -7146 266614
rect -7766 230614 -7146 266058
rect -7766 230058 -7734 230614
rect -7178 230058 -7146 230614
rect -7766 194614 -7146 230058
rect -7766 194058 -7734 194614
rect -7178 194058 -7146 194614
rect -7766 158614 -7146 194058
rect -7766 158058 -7734 158614
rect -7178 158058 -7146 158614
rect -7766 122614 -7146 158058
rect -7766 122058 -7734 122614
rect -7178 122058 -7146 122614
rect -7766 86614 -7146 122058
rect -7766 86058 -7734 86614
rect -7178 86058 -7146 86614
rect -7766 50614 -7146 86058
rect -7766 50058 -7734 50614
rect -7178 50058 -7146 50614
rect -7766 14614 -7146 50058
rect -7766 14058 -7734 14614
rect -7178 14058 -7146 14614
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709082 -6774 709638
rect -6218 709082 -6186 709638
rect -6806 676894 -6186 709082
rect -6806 676338 -6774 676894
rect -6218 676338 -6186 676894
rect -6806 640894 -6186 676338
rect -6806 640338 -6774 640894
rect -6218 640338 -6186 640894
rect -6806 604894 -6186 640338
rect -6806 604338 -6774 604894
rect -6218 604338 -6186 604894
rect -6806 568894 -6186 604338
rect -6806 568338 -6774 568894
rect -6218 568338 -6186 568894
rect -6806 532894 -6186 568338
rect -6806 532338 -6774 532894
rect -6218 532338 -6186 532894
rect -6806 496894 -6186 532338
rect -6806 496338 -6774 496894
rect -6218 496338 -6186 496894
rect -6806 460894 -6186 496338
rect -6806 460338 -6774 460894
rect -6218 460338 -6186 460894
rect -6806 424894 -6186 460338
rect -6806 424338 -6774 424894
rect -6218 424338 -6186 424894
rect -6806 388894 -6186 424338
rect -6806 388338 -6774 388894
rect -6218 388338 -6186 388894
rect -6806 352894 -6186 388338
rect -6806 352338 -6774 352894
rect -6218 352338 -6186 352894
rect -6806 316894 -6186 352338
rect -6806 316338 -6774 316894
rect -6218 316338 -6186 316894
rect -6806 280894 -6186 316338
rect -6806 280338 -6774 280894
rect -6218 280338 -6186 280894
rect -6806 244894 -6186 280338
rect -6806 244338 -6774 244894
rect -6218 244338 -6186 244894
rect -6806 208894 -6186 244338
rect -6806 208338 -6774 208894
rect -6218 208338 -6186 208894
rect -6806 172894 -6186 208338
rect -6806 172338 -6774 172894
rect -6218 172338 -6186 172894
rect -6806 136894 -6186 172338
rect -6806 136338 -6774 136894
rect -6218 136338 -6186 136894
rect -6806 100894 -6186 136338
rect -6806 100338 -6774 100894
rect -6218 100338 -6186 100894
rect -6806 64894 -6186 100338
rect -6806 64338 -6774 64894
rect -6218 64338 -6186 64894
rect -6806 28894 -6186 64338
rect -6806 28338 -6774 28894
rect -6218 28338 -6186 28894
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708122 -5814 708678
rect -5258 708122 -5226 708678
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708122 9266 708678
rect 9822 708122 9854 708678
rect -5846 694338 -5814 694894
rect -5258 694338 -5226 694894
rect -5846 658894 -5226 694338
rect -5846 658338 -5814 658894
rect -5258 658338 -5226 658894
rect -5846 622894 -5226 658338
rect -5846 622338 -5814 622894
rect -5258 622338 -5226 622894
rect -5846 586894 -5226 622338
rect -5846 586338 -5814 586894
rect -5258 586338 -5226 586894
rect -5846 550894 -5226 586338
rect -5846 550338 -5814 550894
rect -5258 550338 -5226 550894
rect -5846 514894 -5226 550338
rect -5846 514338 -5814 514894
rect -5258 514338 -5226 514894
rect -5846 478894 -5226 514338
rect -5846 478338 -5814 478894
rect -5258 478338 -5226 478894
rect -5846 442894 -5226 478338
rect -5846 442338 -5814 442894
rect -5258 442338 -5226 442894
rect -5846 406894 -5226 442338
rect -5846 406338 -5814 406894
rect -5258 406338 -5226 406894
rect -5846 370894 -5226 406338
rect -5846 370338 -5814 370894
rect -5258 370338 -5226 370894
rect -5846 334894 -5226 370338
rect -5846 334338 -5814 334894
rect -5258 334338 -5226 334894
rect -5846 298894 -5226 334338
rect -5846 298338 -5814 298894
rect -5258 298338 -5226 298894
rect -5846 262894 -5226 298338
rect -5846 262338 -5814 262894
rect -5258 262338 -5226 262894
rect -5846 226894 -5226 262338
rect -5846 226338 -5814 226894
rect -5258 226338 -5226 226894
rect -5846 190894 -5226 226338
rect -5846 190338 -5814 190894
rect -5258 190338 -5226 190894
rect -5846 154894 -5226 190338
rect -5846 154338 -5814 154894
rect -5258 154338 -5226 154894
rect -5846 118894 -5226 154338
rect -5846 118338 -5814 118894
rect -5258 118338 -5226 118894
rect -5846 82894 -5226 118338
rect -5846 82338 -5814 82894
rect -5258 82338 -5226 82894
rect -5846 46894 -5226 82338
rect -5846 46338 -5814 46894
rect -5258 46338 -5226 46894
rect -5846 10894 -5226 46338
rect -5846 10338 -5814 10894
rect -5258 10338 -5226 10894
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707162 -4854 707718
rect -4298 707162 -4266 707718
rect -4886 673174 -4266 707162
rect -4886 672618 -4854 673174
rect -4298 672618 -4266 673174
rect -4886 637174 -4266 672618
rect -4886 636618 -4854 637174
rect -4298 636618 -4266 637174
rect -4886 601174 -4266 636618
rect -4886 600618 -4854 601174
rect -4298 600618 -4266 601174
rect -4886 565174 -4266 600618
rect -4886 564618 -4854 565174
rect -4298 564618 -4266 565174
rect -4886 529174 -4266 564618
rect -4886 528618 -4854 529174
rect -4298 528618 -4266 529174
rect -4886 493174 -4266 528618
rect -4886 492618 -4854 493174
rect -4298 492618 -4266 493174
rect -4886 457174 -4266 492618
rect -4886 456618 -4854 457174
rect -4298 456618 -4266 457174
rect -4886 421174 -4266 456618
rect -4886 420618 -4854 421174
rect -4298 420618 -4266 421174
rect -4886 385174 -4266 420618
rect -4886 384618 -4854 385174
rect -4298 384618 -4266 385174
rect -4886 349174 -4266 384618
rect -4886 348618 -4854 349174
rect -4298 348618 -4266 349174
rect -4886 313174 -4266 348618
rect -4886 312618 -4854 313174
rect -4298 312618 -4266 313174
rect -4886 277174 -4266 312618
rect -4886 276618 -4854 277174
rect -4298 276618 -4266 277174
rect -4886 241174 -4266 276618
rect -4886 240618 -4854 241174
rect -4298 240618 -4266 241174
rect -4886 205174 -4266 240618
rect -4886 204618 -4854 205174
rect -4298 204618 -4266 205174
rect -4886 169174 -4266 204618
rect -4886 168618 -4854 169174
rect -4298 168618 -4266 169174
rect -4886 133174 -4266 168618
rect -4886 132618 -4854 133174
rect -4298 132618 -4266 133174
rect -4886 97174 -4266 132618
rect -4886 96618 -4854 97174
rect -4298 96618 -4266 97174
rect -4886 61174 -4266 96618
rect -4886 60618 -4854 61174
rect -4298 60618 -4266 61174
rect -4886 25174 -4266 60618
rect -4886 24618 -4854 25174
rect -4298 24618 -4266 25174
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706202 -3894 706758
rect -3338 706202 -3306 706758
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706202 5546 706758
rect 6102 706202 6134 706758
rect -3926 690618 -3894 691174
rect -3338 690618 -3306 691174
rect -3926 655174 -3306 690618
rect -3926 654618 -3894 655174
rect -3338 654618 -3306 655174
rect -3926 619174 -3306 654618
rect -3926 618618 -3894 619174
rect -3338 618618 -3306 619174
rect -3926 583174 -3306 618618
rect -3926 582618 -3894 583174
rect -3338 582618 -3306 583174
rect -3926 547174 -3306 582618
rect -3926 546618 -3894 547174
rect -3338 546618 -3306 547174
rect -3926 511174 -3306 546618
rect -3926 510618 -3894 511174
rect -3338 510618 -3306 511174
rect -3926 475174 -3306 510618
rect -3926 474618 -3894 475174
rect -3338 474618 -3306 475174
rect -3926 439174 -3306 474618
rect -3926 438618 -3894 439174
rect -3338 438618 -3306 439174
rect -3926 403174 -3306 438618
rect -3926 402618 -3894 403174
rect -3338 402618 -3306 403174
rect -3926 367174 -3306 402618
rect -3926 366618 -3894 367174
rect -3338 366618 -3306 367174
rect -3926 331174 -3306 366618
rect -3926 330618 -3894 331174
rect -3338 330618 -3306 331174
rect -3926 295174 -3306 330618
rect -3926 294618 -3894 295174
rect -3338 294618 -3306 295174
rect -3926 259174 -3306 294618
rect -3926 258618 -3894 259174
rect -3338 258618 -3306 259174
rect -3926 223174 -3306 258618
rect -3926 222618 -3894 223174
rect -3338 222618 -3306 223174
rect -3926 187174 -3306 222618
rect -3926 186618 -3894 187174
rect -3338 186618 -3306 187174
rect -3926 151174 -3306 186618
rect -3926 150618 -3894 151174
rect -3338 150618 -3306 151174
rect -3926 115174 -3306 150618
rect -3926 114618 -3894 115174
rect -3338 114618 -3306 115174
rect -3926 79174 -3306 114618
rect -3926 78618 -3894 79174
rect -3338 78618 -3306 79174
rect -3926 43174 -3306 78618
rect -3926 42618 -3894 43174
rect -3338 42618 -3306 43174
rect -3926 7174 -3306 42618
rect -3926 6618 -3894 7174
rect -3338 6618 -3306 7174
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705242 -2934 705798
rect -2378 705242 -2346 705798
rect -2966 669454 -2346 705242
rect -2966 668898 -2934 669454
rect -2378 668898 -2346 669454
rect -2966 633454 -2346 668898
rect -2966 632898 -2934 633454
rect -2378 632898 -2346 633454
rect -2966 597454 -2346 632898
rect -2966 596898 -2934 597454
rect -2378 596898 -2346 597454
rect -2966 561454 -2346 596898
rect -2966 560898 -2934 561454
rect -2378 560898 -2346 561454
rect -2966 525454 -2346 560898
rect -2966 524898 -2934 525454
rect -2378 524898 -2346 525454
rect -2966 489454 -2346 524898
rect -2966 488898 -2934 489454
rect -2378 488898 -2346 489454
rect -2966 453454 -2346 488898
rect -2966 452898 -2934 453454
rect -2378 452898 -2346 453454
rect -2966 417454 -2346 452898
rect -2966 416898 -2934 417454
rect -2378 416898 -2346 417454
rect -2966 381454 -2346 416898
rect -2966 380898 -2934 381454
rect -2378 380898 -2346 381454
rect -2966 345454 -2346 380898
rect -2966 344898 -2934 345454
rect -2378 344898 -2346 345454
rect -2966 309454 -2346 344898
rect -2966 308898 -2934 309454
rect -2378 308898 -2346 309454
rect -2966 273454 -2346 308898
rect -2966 272898 -2934 273454
rect -2378 272898 -2346 273454
rect -2966 237454 -2346 272898
rect -2966 236898 -2934 237454
rect -2378 236898 -2346 237454
rect -2966 201454 -2346 236898
rect -2966 200898 -2934 201454
rect -2378 200898 -2346 201454
rect -2966 165454 -2346 200898
rect -2966 164898 -2934 165454
rect -2378 164898 -2346 165454
rect -2966 129454 -2346 164898
rect -2966 128898 -2934 129454
rect -2378 128898 -2346 129454
rect -2966 93454 -2346 128898
rect -2966 92898 -2934 93454
rect -2378 92898 -2346 93454
rect -2966 57454 -2346 92898
rect -2966 56898 -2934 57454
rect -2378 56898 -2346 57454
rect -2966 21454 -2346 56898
rect -2966 20898 -2934 21454
rect -2378 20898 -2346 21454
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704282 -1974 704838
rect -1418 704282 -1386 704838
rect -2006 687454 -1386 704282
rect -2006 686898 -1974 687454
rect -1418 686898 -1386 687454
rect -2006 651454 -1386 686898
rect -2006 650898 -1974 651454
rect -1418 650898 -1386 651454
rect -2006 615454 -1386 650898
rect -2006 614898 -1974 615454
rect -1418 614898 -1386 615454
rect -2006 579454 -1386 614898
rect -2006 578898 -1974 579454
rect -1418 578898 -1386 579454
rect -2006 543454 -1386 578898
rect -2006 542898 -1974 543454
rect -1418 542898 -1386 543454
rect -2006 507454 -1386 542898
rect -2006 506898 -1974 507454
rect -1418 506898 -1386 507454
rect -2006 471454 -1386 506898
rect -2006 470898 -1974 471454
rect -1418 470898 -1386 471454
rect -2006 435454 -1386 470898
rect -2006 434898 -1974 435454
rect -1418 434898 -1386 435454
rect -2006 399454 -1386 434898
rect -2006 398898 -1974 399454
rect -1418 398898 -1386 399454
rect -2006 363454 -1386 398898
rect -2006 362898 -1974 363454
rect -1418 362898 -1386 363454
rect -2006 327454 -1386 362898
rect -2006 326898 -1974 327454
rect -1418 326898 -1386 327454
rect -2006 291454 -1386 326898
rect -2006 290898 -1974 291454
rect -1418 290898 -1386 291454
rect -2006 255454 -1386 290898
rect -2006 254898 -1974 255454
rect -1418 254898 -1386 255454
rect -2006 219454 -1386 254898
rect -2006 218898 -1974 219454
rect -1418 218898 -1386 219454
rect -2006 183454 -1386 218898
rect -2006 182898 -1974 183454
rect -1418 182898 -1386 183454
rect -2006 147454 -1386 182898
rect -2006 146898 -1974 147454
rect -1418 146898 -1386 147454
rect -2006 111454 -1386 146898
rect -2006 110898 -1974 111454
rect -1418 110898 -1386 111454
rect -2006 75454 -1386 110898
rect -2006 74898 -1974 75454
rect -1418 74898 -1386 75454
rect -2006 39454 -1386 74898
rect -2006 38898 -1974 39454
rect -1418 38898 -1386 39454
rect -2006 3454 -1386 38898
rect -2006 2898 -1974 3454
rect -1418 2898 -1386 3454
rect -2006 -346 -1386 2898
rect -2006 -902 -1974 -346
rect -1418 -902 -1386 -346
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704282 1826 704838
rect 2382 704282 2414 704838
rect 1794 687454 2414 704282
rect 1794 686898 1826 687454
rect 2382 686898 2414 687454
rect 1794 651454 2414 686898
rect 1794 650898 1826 651454
rect 2382 650898 2414 651454
rect 1794 615454 2414 650898
rect 1794 614898 1826 615454
rect 2382 614898 2414 615454
rect 1794 579454 2414 614898
rect 1794 578898 1826 579454
rect 2382 578898 2414 579454
rect 1794 543454 2414 578898
rect 1794 542898 1826 543454
rect 2382 542898 2414 543454
rect 1794 507454 2414 542898
rect 1794 506898 1826 507454
rect 2382 506898 2414 507454
rect 1794 471454 2414 506898
rect 1794 470898 1826 471454
rect 2382 470898 2414 471454
rect 1794 435454 2414 470898
rect 1794 434898 1826 435454
rect 2382 434898 2414 435454
rect 1794 399454 2414 434898
rect 1794 398898 1826 399454
rect 2382 398898 2414 399454
rect 1794 363454 2414 398898
rect 1794 362898 1826 363454
rect 2382 362898 2414 363454
rect 1794 327454 2414 362898
rect 1794 326898 1826 327454
rect 2382 326898 2414 327454
rect 1794 291454 2414 326898
rect 1794 290898 1826 291454
rect 2382 290898 2414 291454
rect 1794 255454 2414 290898
rect 1794 254898 1826 255454
rect 2382 254898 2414 255454
rect 1794 219454 2414 254898
rect 1794 218898 1826 219454
rect 2382 218898 2414 219454
rect 1794 183454 2414 218898
rect 1794 182898 1826 183454
rect 2382 182898 2414 183454
rect 1794 147454 2414 182898
rect 1794 146898 1826 147454
rect 2382 146898 2414 147454
rect 1794 111454 2414 146898
rect 1794 110898 1826 111454
rect 2382 110898 2414 111454
rect 1794 75454 2414 110898
rect 1794 74898 1826 75454
rect 2382 74898 2414 75454
rect 1794 39454 2414 74898
rect 1794 38898 1826 39454
rect 2382 38898 2414 39454
rect 1794 3454 2414 38898
rect 1794 2898 1826 3454
rect 2382 2898 2414 3454
rect 1794 -346 2414 2898
rect 1794 -902 1826 -346
rect 2382 -902 2414 -346
rect -2966 -1862 -2934 -1306
rect -2378 -1862 -2346 -1306
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690618 5546 691174
rect 6102 690618 6134 691174
rect 5514 655174 6134 690618
rect 5514 654618 5546 655174
rect 6102 654618 6134 655174
rect 5514 619174 6134 654618
rect 5514 618618 5546 619174
rect 6102 618618 6134 619174
rect 5514 583174 6134 618618
rect 5514 582618 5546 583174
rect 6102 582618 6134 583174
rect 5514 547174 6134 582618
rect 5514 546618 5546 547174
rect 6102 546618 6134 547174
rect 5514 511174 6134 546618
rect 5514 510618 5546 511174
rect 6102 510618 6134 511174
rect 5514 475174 6134 510618
rect 5514 474618 5546 475174
rect 6102 474618 6134 475174
rect 5514 439174 6134 474618
rect 5514 438618 5546 439174
rect 6102 438618 6134 439174
rect 5514 403174 6134 438618
rect 5514 402618 5546 403174
rect 6102 402618 6134 403174
rect 5514 367174 6134 402618
rect 5514 366618 5546 367174
rect 6102 366618 6134 367174
rect 5514 331174 6134 366618
rect 5514 330618 5546 331174
rect 6102 330618 6134 331174
rect 5514 295174 6134 330618
rect 5514 294618 5546 295174
rect 6102 294618 6134 295174
rect 5514 259174 6134 294618
rect 5514 258618 5546 259174
rect 6102 258618 6134 259174
rect 5514 223174 6134 258618
rect 5514 222618 5546 223174
rect 6102 222618 6134 223174
rect 5514 187174 6134 222618
rect 5514 186618 5546 187174
rect 6102 186618 6134 187174
rect 5514 151174 6134 186618
rect 5514 150618 5546 151174
rect 6102 150618 6134 151174
rect 5514 115174 6134 150618
rect 5514 114618 5546 115174
rect 6102 114618 6134 115174
rect 5514 79174 6134 114618
rect 5514 78618 5546 79174
rect 6102 78618 6134 79174
rect 5514 43174 6134 78618
rect 5514 42618 5546 43174
rect 6102 42618 6134 43174
rect 5514 7174 6134 42618
rect 5514 6618 5546 7174
rect 6102 6618 6134 7174
rect -3926 -2822 -3894 -2266
rect -3338 -2822 -3306 -2266
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2822 5546 -2266
rect 6102 -2822 6134 -2266
rect -4886 -3782 -4854 -3226
rect -4298 -3782 -4266 -3226
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694338 9266 694894
rect 9822 694338 9854 694894
rect 9234 658894 9854 694338
rect 9234 658338 9266 658894
rect 9822 658338 9854 658894
rect 9234 622894 9854 658338
rect 9234 622338 9266 622894
rect 9822 622338 9854 622894
rect 9234 586894 9854 622338
rect 9234 586338 9266 586894
rect 9822 586338 9854 586894
rect 9234 550894 9854 586338
rect 9234 550338 9266 550894
rect 9822 550338 9854 550894
rect 9234 514894 9854 550338
rect 9234 514338 9266 514894
rect 9822 514338 9854 514894
rect 9234 478894 9854 514338
rect 9234 478338 9266 478894
rect 9822 478338 9854 478894
rect 9234 442894 9854 478338
rect 9234 442338 9266 442894
rect 9822 442338 9854 442894
rect 9234 406894 9854 442338
rect 9234 406338 9266 406894
rect 9822 406338 9854 406894
rect 9234 370894 9854 406338
rect 9234 370338 9266 370894
rect 9822 370338 9854 370894
rect 9234 334894 9854 370338
rect 9234 334338 9266 334894
rect 9822 334338 9854 334894
rect 9234 298894 9854 334338
rect 9234 298338 9266 298894
rect 9822 298338 9854 298894
rect 9234 262894 9854 298338
rect 9234 262338 9266 262894
rect 9822 262338 9854 262894
rect 9234 226894 9854 262338
rect 9234 226338 9266 226894
rect 9822 226338 9854 226894
rect 9234 190894 9854 226338
rect 9234 190338 9266 190894
rect 9822 190338 9854 190894
rect 9234 154894 9854 190338
rect 9234 154338 9266 154894
rect 9822 154338 9854 154894
rect 9234 118894 9854 154338
rect 9234 118338 9266 118894
rect 9822 118338 9854 118894
rect 9234 82894 9854 118338
rect 9234 82338 9266 82894
rect 9822 82338 9854 82894
rect 9234 46894 9854 82338
rect 9234 46338 9266 46894
rect 9822 46338 9854 46894
rect 9234 10894 9854 46338
rect 9234 10338 9266 10894
rect 9822 10338 9854 10894
rect -5846 -4742 -5814 -4186
rect -5258 -4742 -5226 -4186
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4742 9266 -4186
rect 9822 -4742 9854 -4186
rect -6806 -5702 -6774 -5146
rect -6218 -5702 -6186 -5146
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711002 30986 711558
rect 31542 711002 31574 711558
rect 27234 709638 27854 709670
rect 27234 709082 27266 709638
rect 27822 709082 27854 709638
rect 23514 707718 24134 707750
rect 23514 707162 23546 707718
rect 24102 707162 24134 707718
rect 12954 698058 12986 698614
rect 13542 698058 13574 698614
rect 12954 662614 13574 698058
rect 12954 662058 12986 662614
rect 13542 662058 13574 662614
rect 12954 626614 13574 662058
rect 12954 626058 12986 626614
rect 13542 626058 13574 626614
rect 12954 590614 13574 626058
rect 12954 590058 12986 590614
rect 13542 590058 13574 590614
rect 12954 554614 13574 590058
rect 12954 554058 12986 554614
rect 13542 554058 13574 554614
rect 12954 518614 13574 554058
rect 12954 518058 12986 518614
rect 13542 518058 13574 518614
rect 12954 482614 13574 518058
rect 12954 482058 12986 482614
rect 13542 482058 13574 482614
rect 12954 446614 13574 482058
rect 12954 446058 12986 446614
rect 13542 446058 13574 446614
rect 12954 410614 13574 446058
rect 12954 410058 12986 410614
rect 13542 410058 13574 410614
rect 12954 374614 13574 410058
rect 12954 374058 12986 374614
rect 13542 374058 13574 374614
rect 12954 338614 13574 374058
rect 12954 338058 12986 338614
rect 13542 338058 13574 338614
rect 12954 302614 13574 338058
rect 12954 302058 12986 302614
rect 13542 302058 13574 302614
rect 12954 266614 13574 302058
rect 12954 266058 12986 266614
rect 13542 266058 13574 266614
rect 12954 230614 13574 266058
rect 12954 230058 12986 230614
rect 13542 230058 13574 230614
rect 12954 194614 13574 230058
rect 12954 194058 12986 194614
rect 13542 194058 13574 194614
rect 12954 158614 13574 194058
rect 12954 158058 12986 158614
rect 13542 158058 13574 158614
rect 12954 122614 13574 158058
rect 12954 122058 12986 122614
rect 13542 122058 13574 122614
rect 12954 86614 13574 122058
rect 12954 86058 12986 86614
rect 13542 86058 13574 86614
rect 12954 50614 13574 86058
rect 12954 50058 12986 50614
rect 13542 50058 13574 50614
rect 12954 14614 13574 50058
rect 12954 14058 12986 14614
rect 13542 14058 13574 14614
rect -7766 -6662 -7734 -6106
rect -7178 -6662 -7146 -6106
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705242 19826 705798
rect 20382 705242 20414 705798
rect 19794 669454 20414 705242
rect 19794 668898 19826 669454
rect 20382 668898 20414 669454
rect 19794 633454 20414 668898
rect 19794 632898 19826 633454
rect 20382 632898 20414 633454
rect 19794 597454 20414 632898
rect 19794 596898 19826 597454
rect 20382 596898 20414 597454
rect 19794 561454 20414 596898
rect 19794 560898 19826 561454
rect 20382 560898 20414 561454
rect 19794 525454 20414 560898
rect 19794 524898 19826 525454
rect 20382 524898 20414 525454
rect 19794 489454 20414 524898
rect 19794 488898 19826 489454
rect 20382 488898 20414 489454
rect 19794 453454 20414 488898
rect 19794 452898 19826 453454
rect 20382 452898 20414 453454
rect 19794 417454 20414 452898
rect 19794 416898 19826 417454
rect 20382 416898 20414 417454
rect 19794 381454 20414 416898
rect 19794 380898 19826 381454
rect 20382 380898 20414 381454
rect 19794 345454 20414 380898
rect 19794 344898 19826 345454
rect 20382 344898 20414 345454
rect 19794 309454 20414 344898
rect 19794 308898 19826 309454
rect 20382 308898 20414 309454
rect 19794 273454 20414 308898
rect 19794 272898 19826 273454
rect 20382 272898 20414 273454
rect 19794 237454 20414 272898
rect 19794 236898 19826 237454
rect 20382 236898 20414 237454
rect 19794 201454 20414 236898
rect 19794 200898 19826 201454
rect 20382 200898 20414 201454
rect 19794 165454 20414 200898
rect 19794 164898 19826 165454
rect 20382 164898 20414 165454
rect 19794 129454 20414 164898
rect 19794 128898 19826 129454
rect 20382 128898 20414 129454
rect 19794 93454 20414 128898
rect 19794 92898 19826 93454
rect 20382 92898 20414 93454
rect 19794 57454 20414 92898
rect 19794 56898 19826 57454
rect 20382 56898 20414 57454
rect 19794 21454 20414 56898
rect 19794 20898 19826 21454
rect 20382 20898 20414 21454
rect 19794 -1306 20414 20898
rect 19794 -1862 19826 -1306
rect 20382 -1862 20414 -1306
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672618 23546 673174
rect 24102 672618 24134 673174
rect 23514 637174 24134 672618
rect 23514 636618 23546 637174
rect 24102 636618 24134 637174
rect 23514 601174 24134 636618
rect 23514 600618 23546 601174
rect 24102 600618 24134 601174
rect 23514 565174 24134 600618
rect 23514 564618 23546 565174
rect 24102 564618 24134 565174
rect 23514 529174 24134 564618
rect 23514 528618 23546 529174
rect 24102 528618 24134 529174
rect 23514 493174 24134 528618
rect 23514 492618 23546 493174
rect 24102 492618 24134 493174
rect 23514 457174 24134 492618
rect 23514 456618 23546 457174
rect 24102 456618 24134 457174
rect 23514 421174 24134 456618
rect 23514 420618 23546 421174
rect 24102 420618 24134 421174
rect 23514 385174 24134 420618
rect 23514 384618 23546 385174
rect 24102 384618 24134 385174
rect 23514 349174 24134 384618
rect 23514 348618 23546 349174
rect 24102 348618 24134 349174
rect 23514 313174 24134 348618
rect 23514 312618 23546 313174
rect 24102 312618 24134 313174
rect 23514 277174 24134 312618
rect 23514 276618 23546 277174
rect 24102 276618 24134 277174
rect 23514 241174 24134 276618
rect 23514 240618 23546 241174
rect 24102 240618 24134 241174
rect 23514 205174 24134 240618
rect 23514 204618 23546 205174
rect 24102 204618 24134 205174
rect 23514 169174 24134 204618
rect 23514 168618 23546 169174
rect 24102 168618 24134 169174
rect 23514 133174 24134 168618
rect 23514 132618 23546 133174
rect 24102 132618 24134 133174
rect 23514 97174 24134 132618
rect 23514 96618 23546 97174
rect 24102 96618 24134 97174
rect 23514 61174 24134 96618
rect 23514 60618 23546 61174
rect 24102 60618 24134 61174
rect 23514 25174 24134 60618
rect 23514 24618 23546 25174
rect 24102 24618 24134 25174
rect 23514 -3226 24134 24618
rect 23514 -3782 23546 -3226
rect 24102 -3782 24134 -3226
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676338 27266 676894
rect 27822 676338 27854 676894
rect 27234 640894 27854 676338
rect 27234 640338 27266 640894
rect 27822 640338 27854 640894
rect 27234 604894 27854 640338
rect 27234 604338 27266 604894
rect 27822 604338 27854 604894
rect 27234 568894 27854 604338
rect 27234 568338 27266 568894
rect 27822 568338 27854 568894
rect 27234 532894 27854 568338
rect 27234 532338 27266 532894
rect 27822 532338 27854 532894
rect 27234 496894 27854 532338
rect 27234 496338 27266 496894
rect 27822 496338 27854 496894
rect 27234 460894 27854 496338
rect 27234 460338 27266 460894
rect 27822 460338 27854 460894
rect 27234 424894 27854 460338
rect 27234 424338 27266 424894
rect 27822 424338 27854 424894
rect 27234 388894 27854 424338
rect 27234 388338 27266 388894
rect 27822 388338 27854 388894
rect 27234 352894 27854 388338
rect 27234 352338 27266 352894
rect 27822 352338 27854 352894
rect 27234 316894 27854 352338
rect 27234 316338 27266 316894
rect 27822 316338 27854 316894
rect 27234 280894 27854 316338
rect 27234 280338 27266 280894
rect 27822 280338 27854 280894
rect 27234 244894 27854 280338
rect 27234 244338 27266 244894
rect 27822 244338 27854 244894
rect 27234 208894 27854 244338
rect 27234 208338 27266 208894
rect 27822 208338 27854 208894
rect 27234 172894 27854 208338
rect 27234 172338 27266 172894
rect 27822 172338 27854 172894
rect 27234 136894 27854 172338
rect 27234 136338 27266 136894
rect 27822 136338 27854 136894
rect 27234 100894 27854 136338
rect 27234 100338 27266 100894
rect 27822 100338 27854 100894
rect 27234 64894 27854 100338
rect 27234 64338 27266 64894
rect 27822 64338 27854 64894
rect 27234 28894 27854 64338
rect 27234 28338 27266 28894
rect 27822 28338 27854 28894
rect 27234 -5146 27854 28338
rect 27234 -5702 27266 -5146
rect 27822 -5702 27854 -5146
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710042 48986 710598
rect 49542 710042 49574 710598
rect 45234 708678 45854 709670
rect 45234 708122 45266 708678
rect 45822 708122 45854 708678
rect 41514 706758 42134 707750
rect 41514 706202 41546 706758
rect 42102 706202 42134 706758
rect 30954 680058 30986 680614
rect 31542 680058 31574 680614
rect 30954 644614 31574 680058
rect 30954 644058 30986 644614
rect 31542 644058 31574 644614
rect 30954 608614 31574 644058
rect 30954 608058 30986 608614
rect 31542 608058 31574 608614
rect 30954 572614 31574 608058
rect 30954 572058 30986 572614
rect 31542 572058 31574 572614
rect 30954 536614 31574 572058
rect 30954 536058 30986 536614
rect 31542 536058 31574 536614
rect 30954 500614 31574 536058
rect 30954 500058 30986 500614
rect 31542 500058 31574 500614
rect 30954 464614 31574 500058
rect 30954 464058 30986 464614
rect 31542 464058 31574 464614
rect 30954 428614 31574 464058
rect 30954 428058 30986 428614
rect 31542 428058 31574 428614
rect 30954 392614 31574 428058
rect 30954 392058 30986 392614
rect 31542 392058 31574 392614
rect 30954 356614 31574 392058
rect 30954 356058 30986 356614
rect 31542 356058 31574 356614
rect 30954 320614 31574 356058
rect 30954 320058 30986 320614
rect 31542 320058 31574 320614
rect 30954 284614 31574 320058
rect 30954 284058 30986 284614
rect 31542 284058 31574 284614
rect 30954 248614 31574 284058
rect 30954 248058 30986 248614
rect 31542 248058 31574 248614
rect 30954 212614 31574 248058
rect 30954 212058 30986 212614
rect 31542 212058 31574 212614
rect 30954 176614 31574 212058
rect 30954 176058 30986 176614
rect 31542 176058 31574 176614
rect 30954 140614 31574 176058
rect 30954 140058 30986 140614
rect 31542 140058 31574 140614
rect 30954 104614 31574 140058
rect 30954 104058 30986 104614
rect 31542 104058 31574 104614
rect 30954 68614 31574 104058
rect 30954 68058 30986 68614
rect 31542 68058 31574 68614
rect 30954 32614 31574 68058
rect 30954 32058 30986 32614
rect 31542 32058 31574 32614
rect 12954 -6662 12986 -6106
rect 13542 -6662 13574 -6106
rect -8726 -7622 -8694 -7066
rect -8138 -7622 -8106 -7066
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704282 37826 704838
rect 38382 704282 38414 704838
rect 37794 687454 38414 704282
rect 37794 686898 37826 687454
rect 38382 686898 38414 687454
rect 37794 651454 38414 686898
rect 37794 650898 37826 651454
rect 38382 650898 38414 651454
rect 37794 615454 38414 650898
rect 37794 614898 37826 615454
rect 38382 614898 38414 615454
rect 37794 579454 38414 614898
rect 37794 578898 37826 579454
rect 38382 578898 38414 579454
rect 37794 543454 38414 578898
rect 37794 542898 37826 543454
rect 38382 542898 38414 543454
rect 37794 507454 38414 542898
rect 37794 506898 37826 507454
rect 38382 506898 38414 507454
rect 37794 471454 38414 506898
rect 37794 470898 37826 471454
rect 38382 470898 38414 471454
rect 37794 435454 38414 470898
rect 37794 434898 37826 435454
rect 38382 434898 38414 435454
rect 37794 399454 38414 434898
rect 37794 398898 37826 399454
rect 38382 398898 38414 399454
rect 37794 363454 38414 398898
rect 37794 362898 37826 363454
rect 38382 362898 38414 363454
rect 37794 327454 38414 362898
rect 37794 326898 37826 327454
rect 38382 326898 38414 327454
rect 37794 291454 38414 326898
rect 37794 290898 37826 291454
rect 38382 290898 38414 291454
rect 37794 255454 38414 290898
rect 37794 254898 37826 255454
rect 38382 254898 38414 255454
rect 37794 219454 38414 254898
rect 37794 218898 37826 219454
rect 38382 218898 38414 219454
rect 37794 183454 38414 218898
rect 37794 182898 37826 183454
rect 38382 182898 38414 183454
rect 37794 147454 38414 182898
rect 37794 146898 37826 147454
rect 38382 146898 38414 147454
rect 37794 111454 38414 146898
rect 37794 110898 37826 111454
rect 38382 110898 38414 111454
rect 37794 75454 38414 110898
rect 37794 74898 37826 75454
rect 38382 74898 38414 75454
rect 37794 39454 38414 74898
rect 37794 38898 37826 39454
rect 38382 38898 38414 39454
rect 37794 3454 38414 38898
rect 37794 2898 37826 3454
rect 38382 2898 38414 3454
rect 37794 -346 38414 2898
rect 37794 -902 37826 -346
rect 38382 -902 38414 -346
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690618 41546 691174
rect 42102 690618 42134 691174
rect 41514 655174 42134 690618
rect 41514 654618 41546 655174
rect 42102 654618 42134 655174
rect 41514 619174 42134 654618
rect 41514 618618 41546 619174
rect 42102 618618 42134 619174
rect 41514 583174 42134 618618
rect 41514 582618 41546 583174
rect 42102 582618 42134 583174
rect 41514 547174 42134 582618
rect 41514 546618 41546 547174
rect 42102 546618 42134 547174
rect 41514 511174 42134 546618
rect 41514 510618 41546 511174
rect 42102 510618 42134 511174
rect 41514 475174 42134 510618
rect 41514 474618 41546 475174
rect 42102 474618 42134 475174
rect 41514 439174 42134 474618
rect 41514 438618 41546 439174
rect 42102 438618 42134 439174
rect 41514 403174 42134 438618
rect 41514 402618 41546 403174
rect 42102 402618 42134 403174
rect 41514 367174 42134 402618
rect 41514 366618 41546 367174
rect 42102 366618 42134 367174
rect 41514 331174 42134 366618
rect 41514 330618 41546 331174
rect 42102 330618 42134 331174
rect 41514 295174 42134 330618
rect 41514 294618 41546 295174
rect 42102 294618 42134 295174
rect 41514 259174 42134 294618
rect 41514 258618 41546 259174
rect 42102 258618 42134 259174
rect 41514 223174 42134 258618
rect 41514 222618 41546 223174
rect 42102 222618 42134 223174
rect 41514 187174 42134 222618
rect 41514 186618 41546 187174
rect 42102 186618 42134 187174
rect 41514 151174 42134 186618
rect 41514 150618 41546 151174
rect 42102 150618 42134 151174
rect 41514 115174 42134 150618
rect 41514 114618 41546 115174
rect 42102 114618 42134 115174
rect 41514 79174 42134 114618
rect 41514 78618 41546 79174
rect 42102 78618 42134 79174
rect 41514 43174 42134 78618
rect 41514 42618 41546 43174
rect 42102 42618 42134 43174
rect 41514 7174 42134 42618
rect 41514 6618 41546 7174
rect 42102 6618 42134 7174
rect 41514 -2266 42134 6618
rect 41514 -2822 41546 -2266
rect 42102 -2822 42134 -2266
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694338 45266 694894
rect 45822 694338 45854 694894
rect 45234 658894 45854 694338
rect 45234 658338 45266 658894
rect 45822 658338 45854 658894
rect 45234 622894 45854 658338
rect 45234 622338 45266 622894
rect 45822 622338 45854 622894
rect 45234 586894 45854 622338
rect 45234 586338 45266 586894
rect 45822 586338 45854 586894
rect 45234 550894 45854 586338
rect 45234 550338 45266 550894
rect 45822 550338 45854 550894
rect 45234 514894 45854 550338
rect 45234 514338 45266 514894
rect 45822 514338 45854 514894
rect 45234 478894 45854 514338
rect 45234 478338 45266 478894
rect 45822 478338 45854 478894
rect 45234 442894 45854 478338
rect 45234 442338 45266 442894
rect 45822 442338 45854 442894
rect 45234 406894 45854 442338
rect 45234 406338 45266 406894
rect 45822 406338 45854 406894
rect 45234 370894 45854 406338
rect 45234 370338 45266 370894
rect 45822 370338 45854 370894
rect 45234 334894 45854 370338
rect 45234 334338 45266 334894
rect 45822 334338 45854 334894
rect 45234 298894 45854 334338
rect 45234 298338 45266 298894
rect 45822 298338 45854 298894
rect 45234 262894 45854 298338
rect 45234 262338 45266 262894
rect 45822 262338 45854 262894
rect 45234 226894 45854 262338
rect 45234 226338 45266 226894
rect 45822 226338 45854 226894
rect 45234 190894 45854 226338
rect 45234 190338 45266 190894
rect 45822 190338 45854 190894
rect 45234 154894 45854 190338
rect 45234 154338 45266 154894
rect 45822 154338 45854 154894
rect 45234 118894 45854 154338
rect 45234 118338 45266 118894
rect 45822 118338 45854 118894
rect 45234 82894 45854 118338
rect 45234 82338 45266 82894
rect 45822 82338 45854 82894
rect 45234 46894 45854 82338
rect 45234 46338 45266 46894
rect 45822 46338 45854 46894
rect 45234 10894 45854 46338
rect 45234 10338 45266 10894
rect 45822 10338 45854 10894
rect 45234 -4186 45854 10338
rect 45234 -4742 45266 -4186
rect 45822 -4742 45854 -4186
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711002 66986 711558
rect 67542 711002 67574 711558
rect 63234 709638 63854 709670
rect 63234 709082 63266 709638
rect 63822 709082 63854 709638
rect 59514 707718 60134 707750
rect 59514 707162 59546 707718
rect 60102 707162 60134 707718
rect 48954 698058 48986 698614
rect 49542 698058 49574 698614
rect 48954 662614 49574 698058
rect 48954 662058 48986 662614
rect 49542 662058 49574 662614
rect 48954 626614 49574 662058
rect 48954 626058 48986 626614
rect 49542 626058 49574 626614
rect 48954 590614 49574 626058
rect 48954 590058 48986 590614
rect 49542 590058 49574 590614
rect 48954 554614 49574 590058
rect 48954 554058 48986 554614
rect 49542 554058 49574 554614
rect 48954 518614 49574 554058
rect 48954 518058 48986 518614
rect 49542 518058 49574 518614
rect 48954 482614 49574 518058
rect 48954 482058 48986 482614
rect 49542 482058 49574 482614
rect 48954 446614 49574 482058
rect 48954 446058 48986 446614
rect 49542 446058 49574 446614
rect 48954 410614 49574 446058
rect 48954 410058 48986 410614
rect 49542 410058 49574 410614
rect 48954 374614 49574 410058
rect 48954 374058 48986 374614
rect 49542 374058 49574 374614
rect 48954 338614 49574 374058
rect 48954 338058 48986 338614
rect 49542 338058 49574 338614
rect 48954 302614 49574 338058
rect 48954 302058 48986 302614
rect 49542 302058 49574 302614
rect 48954 266614 49574 302058
rect 48954 266058 48986 266614
rect 49542 266058 49574 266614
rect 48954 230614 49574 266058
rect 48954 230058 48986 230614
rect 49542 230058 49574 230614
rect 48954 194614 49574 230058
rect 48954 194058 48986 194614
rect 49542 194058 49574 194614
rect 48954 158614 49574 194058
rect 48954 158058 48986 158614
rect 49542 158058 49574 158614
rect 48954 122614 49574 158058
rect 48954 122058 48986 122614
rect 49542 122058 49574 122614
rect 48954 86614 49574 122058
rect 48954 86058 48986 86614
rect 49542 86058 49574 86614
rect 48954 50614 49574 86058
rect 48954 50058 48986 50614
rect 49542 50058 49574 50614
rect 48954 14614 49574 50058
rect 48954 14058 48986 14614
rect 49542 14058 49574 14614
rect 30954 -7622 30986 -7066
rect 31542 -7622 31574 -7066
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705242 55826 705798
rect 56382 705242 56414 705798
rect 55794 669454 56414 705242
rect 55794 668898 55826 669454
rect 56382 668898 56414 669454
rect 55794 633454 56414 668898
rect 55794 632898 55826 633454
rect 56382 632898 56414 633454
rect 55794 597454 56414 632898
rect 55794 596898 55826 597454
rect 56382 596898 56414 597454
rect 55794 561454 56414 596898
rect 55794 560898 55826 561454
rect 56382 560898 56414 561454
rect 55794 525454 56414 560898
rect 55794 524898 55826 525454
rect 56382 524898 56414 525454
rect 55794 489454 56414 524898
rect 55794 488898 55826 489454
rect 56382 488898 56414 489454
rect 55794 453454 56414 488898
rect 55794 452898 55826 453454
rect 56382 452898 56414 453454
rect 55794 417454 56414 452898
rect 55794 416898 55826 417454
rect 56382 416898 56414 417454
rect 55794 381454 56414 416898
rect 55794 380898 55826 381454
rect 56382 380898 56414 381454
rect 55794 345454 56414 380898
rect 55794 344898 55826 345454
rect 56382 344898 56414 345454
rect 55794 309454 56414 344898
rect 55794 308898 55826 309454
rect 56382 308898 56414 309454
rect 55794 273454 56414 308898
rect 55794 272898 55826 273454
rect 56382 272898 56414 273454
rect 55794 237454 56414 272898
rect 55794 236898 55826 237454
rect 56382 236898 56414 237454
rect 55794 201454 56414 236898
rect 55794 200898 55826 201454
rect 56382 200898 56414 201454
rect 55794 165454 56414 200898
rect 55794 164898 55826 165454
rect 56382 164898 56414 165454
rect 55794 129454 56414 164898
rect 55794 128898 55826 129454
rect 56382 128898 56414 129454
rect 55794 93454 56414 128898
rect 55794 92898 55826 93454
rect 56382 92898 56414 93454
rect 55794 57454 56414 92898
rect 55794 56898 55826 57454
rect 56382 56898 56414 57454
rect 55794 21454 56414 56898
rect 55794 20898 55826 21454
rect 56382 20898 56414 21454
rect 55794 -1306 56414 20898
rect 55794 -1862 55826 -1306
rect 56382 -1862 56414 -1306
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672618 59546 673174
rect 60102 672618 60134 673174
rect 59514 637174 60134 672618
rect 59514 636618 59546 637174
rect 60102 636618 60134 637174
rect 59514 601174 60134 636618
rect 59514 600618 59546 601174
rect 60102 600618 60134 601174
rect 59514 565174 60134 600618
rect 59514 564618 59546 565174
rect 60102 564618 60134 565174
rect 59514 529174 60134 564618
rect 59514 528618 59546 529174
rect 60102 528618 60134 529174
rect 59514 493174 60134 528618
rect 59514 492618 59546 493174
rect 60102 492618 60134 493174
rect 59514 457174 60134 492618
rect 59514 456618 59546 457174
rect 60102 456618 60134 457174
rect 59514 421174 60134 456618
rect 59514 420618 59546 421174
rect 60102 420618 60134 421174
rect 59514 385174 60134 420618
rect 59514 384618 59546 385174
rect 60102 384618 60134 385174
rect 59514 349174 60134 384618
rect 59514 348618 59546 349174
rect 60102 348618 60134 349174
rect 59514 313174 60134 348618
rect 59514 312618 59546 313174
rect 60102 312618 60134 313174
rect 59514 277174 60134 312618
rect 59514 276618 59546 277174
rect 60102 276618 60134 277174
rect 59514 241174 60134 276618
rect 59514 240618 59546 241174
rect 60102 240618 60134 241174
rect 59514 205174 60134 240618
rect 59514 204618 59546 205174
rect 60102 204618 60134 205174
rect 59514 169174 60134 204618
rect 59514 168618 59546 169174
rect 60102 168618 60134 169174
rect 59514 133174 60134 168618
rect 59514 132618 59546 133174
rect 60102 132618 60134 133174
rect 59514 97174 60134 132618
rect 59514 96618 59546 97174
rect 60102 96618 60134 97174
rect 59514 61174 60134 96618
rect 59514 60618 59546 61174
rect 60102 60618 60134 61174
rect 59514 25174 60134 60618
rect 59514 24618 59546 25174
rect 60102 24618 60134 25174
rect 59514 -3226 60134 24618
rect 59514 -3782 59546 -3226
rect 60102 -3782 60134 -3226
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676338 63266 676894
rect 63822 676338 63854 676894
rect 63234 640894 63854 676338
rect 63234 640338 63266 640894
rect 63822 640338 63854 640894
rect 63234 604894 63854 640338
rect 63234 604338 63266 604894
rect 63822 604338 63854 604894
rect 63234 568894 63854 604338
rect 63234 568338 63266 568894
rect 63822 568338 63854 568894
rect 63234 532894 63854 568338
rect 63234 532338 63266 532894
rect 63822 532338 63854 532894
rect 63234 496894 63854 532338
rect 63234 496338 63266 496894
rect 63822 496338 63854 496894
rect 63234 460894 63854 496338
rect 63234 460338 63266 460894
rect 63822 460338 63854 460894
rect 63234 424894 63854 460338
rect 63234 424338 63266 424894
rect 63822 424338 63854 424894
rect 63234 388894 63854 424338
rect 63234 388338 63266 388894
rect 63822 388338 63854 388894
rect 63234 352894 63854 388338
rect 63234 352338 63266 352894
rect 63822 352338 63854 352894
rect 63234 316894 63854 352338
rect 63234 316338 63266 316894
rect 63822 316338 63854 316894
rect 63234 280894 63854 316338
rect 63234 280338 63266 280894
rect 63822 280338 63854 280894
rect 63234 244894 63854 280338
rect 63234 244338 63266 244894
rect 63822 244338 63854 244894
rect 63234 208894 63854 244338
rect 63234 208338 63266 208894
rect 63822 208338 63854 208894
rect 63234 172894 63854 208338
rect 63234 172338 63266 172894
rect 63822 172338 63854 172894
rect 63234 136894 63854 172338
rect 63234 136338 63266 136894
rect 63822 136338 63854 136894
rect 63234 100894 63854 136338
rect 63234 100338 63266 100894
rect 63822 100338 63854 100894
rect 63234 64894 63854 100338
rect 63234 64338 63266 64894
rect 63822 64338 63854 64894
rect 63234 28894 63854 64338
rect 63234 28338 63266 28894
rect 63822 28338 63854 28894
rect 63234 -5146 63854 28338
rect 63234 -5702 63266 -5146
rect 63822 -5702 63854 -5146
rect 63234 -5734 63854 -5702
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710042 84986 710598
rect 85542 710042 85574 710598
rect 81234 708678 81854 709670
rect 81234 708122 81266 708678
rect 81822 708122 81854 708678
rect 77514 706758 78134 707750
rect 77514 706202 77546 706758
rect 78102 706202 78134 706758
rect 66954 680058 66986 680614
rect 67542 680058 67574 680614
rect 66954 644614 67574 680058
rect 66954 644058 66986 644614
rect 67542 644058 67574 644614
rect 66954 608614 67574 644058
rect 66954 608058 66986 608614
rect 67542 608058 67574 608614
rect 66954 572614 67574 608058
rect 66954 572058 66986 572614
rect 67542 572058 67574 572614
rect 66954 536614 67574 572058
rect 66954 536058 66986 536614
rect 67542 536058 67574 536614
rect 66954 500614 67574 536058
rect 66954 500058 66986 500614
rect 67542 500058 67574 500614
rect 66954 464614 67574 500058
rect 66954 464058 66986 464614
rect 67542 464058 67574 464614
rect 66954 428614 67574 464058
rect 66954 428058 66986 428614
rect 67542 428058 67574 428614
rect 66954 392614 67574 428058
rect 66954 392058 66986 392614
rect 67542 392058 67574 392614
rect 66954 356614 67574 392058
rect 66954 356058 66986 356614
rect 67542 356058 67574 356614
rect 66954 320614 67574 356058
rect 66954 320058 66986 320614
rect 67542 320058 67574 320614
rect 66954 284614 67574 320058
rect 66954 284058 66986 284614
rect 67542 284058 67574 284614
rect 66954 248614 67574 284058
rect 66954 248058 66986 248614
rect 67542 248058 67574 248614
rect 66954 212614 67574 248058
rect 66954 212058 66986 212614
rect 67542 212058 67574 212614
rect 66954 176614 67574 212058
rect 66954 176058 66986 176614
rect 67542 176058 67574 176614
rect 66954 140614 67574 176058
rect 66954 140058 66986 140614
rect 67542 140058 67574 140614
rect 66954 104614 67574 140058
rect 66954 104058 66986 104614
rect 67542 104058 67574 104614
rect 66954 68614 67574 104058
rect 66954 68058 66986 68614
rect 67542 68058 67574 68614
rect 66954 32614 67574 68058
rect 66954 32058 66986 32614
rect 67542 32058 67574 32614
rect 48954 -6662 48986 -6106
rect 49542 -6662 49574 -6106
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 704838 74414 705830
rect 73794 704282 73826 704838
rect 74382 704282 74414 704838
rect 73794 687454 74414 704282
rect 73794 686898 73826 687454
rect 74382 686898 74414 687454
rect 73794 651454 74414 686898
rect 73794 650898 73826 651454
rect 74382 650898 74414 651454
rect 73794 615454 74414 650898
rect 73794 614898 73826 615454
rect 74382 614898 74414 615454
rect 73794 579454 74414 614898
rect 73794 578898 73826 579454
rect 74382 578898 74414 579454
rect 73794 543454 74414 578898
rect 73794 542898 73826 543454
rect 74382 542898 74414 543454
rect 73794 507454 74414 542898
rect 73794 506898 73826 507454
rect 74382 506898 74414 507454
rect 73794 471454 74414 506898
rect 73794 470898 73826 471454
rect 74382 470898 74414 471454
rect 73794 435454 74414 470898
rect 73794 434898 73826 435454
rect 74382 434898 74414 435454
rect 73794 399454 74414 434898
rect 73794 398898 73826 399454
rect 74382 398898 74414 399454
rect 73794 363454 74414 398898
rect 73794 362898 73826 363454
rect 74382 362898 74414 363454
rect 73794 327454 74414 362898
rect 73794 326898 73826 327454
rect 74382 326898 74414 327454
rect 73794 291454 74414 326898
rect 73794 290898 73826 291454
rect 74382 290898 74414 291454
rect 73794 255454 74414 290898
rect 73794 254898 73826 255454
rect 74382 254898 74414 255454
rect 73794 219454 74414 254898
rect 73794 218898 73826 219454
rect 74382 218898 74414 219454
rect 73794 183454 74414 218898
rect 73794 182898 73826 183454
rect 74382 182898 74414 183454
rect 73794 147454 74414 182898
rect 73794 146898 73826 147454
rect 74382 146898 74414 147454
rect 73794 111454 74414 146898
rect 73794 110898 73826 111454
rect 74382 110898 74414 111454
rect 73794 75454 74414 110898
rect 73794 74898 73826 75454
rect 74382 74898 74414 75454
rect 73794 39454 74414 74898
rect 73794 38898 73826 39454
rect 74382 38898 74414 39454
rect 73794 3454 74414 38898
rect 73794 2898 73826 3454
rect 74382 2898 74414 3454
rect 73794 -346 74414 2898
rect 73794 -902 73826 -346
rect 74382 -902 74414 -346
rect 73794 -1894 74414 -902
rect 77514 691174 78134 706202
rect 77514 690618 77546 691174
rect 78102 690618 78134 691174
rect 77514 655174 78134 690618
rect 77514 654618 77546 655174
rect 78102 654618 78134 655174
rect 77514 619174 78134 654618
rect 77514 618618 77546 619174
rect 78102 618618 78134 619174
rect 77514 583174 78134 618618
rect 77514 582618 77546 583174
rect 78102 582618 78134 583174
rect 77514 547174 78134 582618
rect 77514 546618 77546 547174
rect 78102 546618 78134 547174
rect 77514 511174 78134 546618
rect 77514 510618 77546 511174
rect 78102 510618 78134 511174
rect 77514 475174 78134 510618
rect 77514 474618 77546 475174
rect 78102 474618 78134 475174
rect 77514 439174 78134 474618
rect 77514 438618 77546 439174
rect 78102 438618 78134 439174
rect 77514 403174 78134 438618
rect 77514 402618 77546 403174
rect 78102 402618 78134 403174
rect 77514 367174 78134 402618
rect 77514 366618 77546 367174
rect 78102 366618 78134 367174
rect 77514 331174 78134 366618
rect 77514 330618 77546 331174
rect 78102 330618 78134 331174
rect 77514 295174 78134 330618
rect 77514 294618 77546 295174
rect 78102 294618 78134 295174
rect 77514 259174 78134 294618
rect 77514 258618 77546 259174
rect 78102 258618 78134 259174
rect 77514 223174 78134 258618
rect 77514 222618 77546 223174
rect 78102 222618 78134 223174
rect 77514 187174 78134 222618
rect 77514 186618 77546 187174
rect 78102 186618 78134 187174
rect 77514 151174 78134 186618
rect 77514 150618 77546 151174
rect 78102 150618 78134 151174
rect 77514 115174 78134 150618
rect 77514 114618 77546 115174
rect 78102 114618 78134 115174
rect 77514 79174 78134 114618
rect 77514 78618 77546 79174
rect 78102 78618 78134 79174
rect 77514 43174 78134 78618
rect 77514 42618 77546 43174
rect 78102 42618 78134 43174
rect 77514 7174 78134 42618
rect 77514 6618 77546 7174
rect 78102 6618 78134 7174
rect 77514 -2266 78134 6618
rect 77514 -2822 77546 -2266
rect 78102 -2822 78134 -2266
rect 77514 -3814 78134 -2822
rect 81234 694894 81854 708122
rect 81234 694338 81266 694894
rect 81822 694338 81854 694894
rect 81234 658894 81854 694338
rect 81234 658338 81266 658894
rect 81822 658338 81854 658894
rect 81234 622894 81854 658338
rect 81234 622338 81266 622894
rect 81822 622338 81854 622894
rect 81234 586894 81854 622338
rect 81234 586338 81266 586894
rect 81822 586338 81854 586894
rect 81234 550894 81854 586338
rect 81234 550338 81266 550894
rect 81822 550338 81854 550894
rect 81234 514894 81854 550338
rect 81234 514338 81266 514894
rect 81822 514338 81854 514894
rect 81234 478894 81854 514338
rect 81234 478338 81266 478894
rect 81822 478338 81854 478894
rect 81234 442894 81854 478338
rect 81234 442338 81266 442894
rect 81822 442338 81854 442894
rect 81234 406894 81854 442338
rect 81234 406338 81266 406894
rect 81822 406338 81854 406894
rect 81234 370894 81854 406338
rect 81234 370338 81266 370894
rect 81822 370338 81854 370894
rect 81234 334894 81854 370338
rect 81234 334338 81266 334894
rect 81822 334338 81854 334894
rect 81234 298894 81854 334338
rect 81234 298338 81266 298894
rect 81822 298338 81854 298894
rect 81234 262894 81854 298338
rect 81234 262338 81266 262894
rect 81822 262338 81854 262894
rect 81234 226894 81854 262338
rect 81234 226338 81266 226894
rect 81822 226338 81854 226894
rect 81234 190894 81854 226338
rect 81234 190338 81266 190894
rect 81822 190338 81854 190894
rect 81234 154894 81854 190338
rect 81234 154338 81266 154894
rect 81822 154338 81854 154894
rect 81234 118894 81854 154338
rect 81234 118338 81266 118894
rect 81822 118338 81854 118894
rect 81234 82894 81854 118338
rect 81234 82338 81266 82894
rect 81822 82338 81854 82894
rect 81234 46894 81854 82338
rect 81234 46338 81266 46894
rect 81822 46338 81854 46894
rect 81234 10894 81854 46338
rect 81234 10338 81266 10894
rect 81822 10338 81854 10894
rect 81234 -4186 81854 10338
rect 81234 -4742 81266 -4186
rect 81822 -4742 81854 -4186
rect 81234 -5734 81854 -4742
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711002 102986 711558
rect 103542 711002 103574 711558
rect 99234 709638 99854 709670
rect 99234 709082 99266 709638
rect 99822 709082 99854 709638
rect 95514 707718 96134 707750
rect 95514 707162 95546 707718
rect 96102 707162 96134 707718
rect 84954 698058 84986 698614
rect 85542 698058 85574 698614
rect 84954 662614 85574 698058
rect 84954 662058 84986 662614
rect 85542 662058 85574 662614
rect 84954 626614 85574 662058
rect 84954 626058 84986 626614
rect 85542 626058 85574 626614
rect 84954 590614 85574 626058
rect 84954 590058 84986 590614
rect 85542 590058 85574 590614
rect 84954 554614 85574 590058
rect 84954 554058 84986 554614
rect 85542 554058 85574 554614
rect 84954 518614 85574 554058
rect 84954 518058 84986 518614
rect 85542 518058 85574 518614
rect 84954 482614 85574 518058
rect 84954 482058 84986 482614
rect 85542 482058 85574 482614
rect 84954 446614 85574 482058
rect 84954 446058 84986 446614
rect 85542 446058 85574 446614
rect 84954 410614 85574 446058
rect 84954 410058 84986 410614
rect 85542 410058 85574 410614
rect 84954 374614 85574 410058
rect 84954 374058 84986 374614
rect 85542 374058 85574 374614
rect 84954 338614 85574 374058
rect 84954 338058 84986 338614
rect 85542 338058 85574 338614
rect 84954 302614 85574 338058
rect 84954 302058 84986 302614
rect 85542 302058 85574 302614
rect 84954 266614 85574 302058
rect 84954 266058 84986 266614
rect 85542 266058 85574 266614
rect 84954 230614 85574 266058
rect 84954 230058 84986 230614
rect 85542 230058 85574 230614
rect 84954 194614 85574 230058
rect 84954 194058 84986 194614
rect 85542 194058 85574 194614
rect 84954 158614 85574 194058
rect 84954 158058 84986 158614
rect 85542 158058 85574 158614
rect 84954 122614 85574 158058
rect 84954 122058 84986 122614
rect 85542 122058 85574 122614
rect 84954 86614 85574 122058
rect 84954 86058 84986 86614
rect 85542 86058 85574 86614
rect 84954 50614 85574 86058
rect 84954 50058 84986 50614
rect 85542 50058 85574 50614
rect 84954 14614 85574 50058
rect 84954 14058 84986 14614
rect 85542 14058 85574 14614
rect 66954 -7622 66986 -7066
rect 67542 -7622 67574 -7066
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 705798 92414 705830
rect 91794 705242 91826 705798
rect 92382 705242 92414 705798
rect 91794 669454 92414 705242
rect 91794 668898 91826 669454
rect 92382 668898 92414 669454
rect 91794 633454 92414 668898
rect 91794 632898 91826 633454
rect 92382 632898 92414 633454
rect 91794 597454 92414 632898
rect 91794 596898 91826 597454
rect 92382 596898 92414 597454
rect 91794 561454 92414 596898
rect 91794 560898 91826 561454
rect 92382 560898 92414 561454
rect 91794 525454 92414 560898
rect 91794 524898 91826 525454
rect 92382 524898 92414 525454
rect 91794 489454 92414 524898
rect 91794 488898 91826 489454
rect 92382 488898 92414 489454
rect 91794 453454 92414 488898
rect 91794 452898 91826 453454
rect 92382 452898 92414 453454
rect 91794 417454 92414 452898
rect 91794 416898 91826 417454
rect 92382 416898 92414 417454
rect 91794 381454 92414 416898
rect 91794 380898 91826 381454
rect 92382 380898 92414 381454
rect 91794 345454 92414 380898
rect 91794 344898 91826 345454
rect 92382 344898 92414 345454
rect 91794 309454 92414 344898
rect 91794 308898 91826 309454
rect 92382 308898 92414 309454
rect 91794 273454 92414 308898
rect 91794 272898 91826 273454
rect 92382 272898 92414 273454
rect 91794 237454 92414 272898
rect 91794 236898 91826 237454
rect 92382 236898 92414 237454
rect 91794 201454 92414 236898
rect 91794 200898 91826 201454
rect 92382 200898 92414 201454
rect 91794 165454 92414 200898
rect 91794 164898 91826 165454
rect 92382 164898 92414 165454
rect 91794 129454 92414 164898
rect 91794 128898 91826 129454
rect 92382 128898 92414 129454
rect 91794 93454 92414 128898
rect 91794 92898 91826 93454
rect 92382 92898 92414 93454
rect 91794 57454 92414 92898
rect 91794 56898 91826 57454
rect 92382 56898 92414 57454
rect 91794 21454 92414 56898
rect 91794 20898 91826 21454
rect 92382 20898 92414 21454
rect 91794 -1306 92414 20898
rect 91794 -1862 91826 -1306
rect 92382 -1862 92414 -1306
rect 91794 -1894 92414 -1862
rect 95514 673174 96134 707162
rect 95514 672618 95546 673174
rect 96102 672618 96134 673174
rect 95514 637174 96134 672618
rect 95514 636618 95546 637174
rect 96102 636618 96134 637174
rect 95514 601174 96134 636618
rect 95514 600618 95546 601174
rect 96102 600618 96134 601174
rect 95514 565174 96134 600618
rect 95514 564618 95546 565174
rect 96102 564618 96134 565174
rect 95514 529174 96134 564618
rect 95514 528618 95546 529174
rect 96102 528618 96134 529174
rect 95514 493174 96134 528618
rect 95514 492618 95546 493174
rect 96102 492618 96134 493174
rect 95514 457174 96134 492618
rect 95514 456618 95546 457174
rect 96102 456618 96134 457174
rect 95514 421174 96134 456618
rect 95514 420618 95546 421174
rect 96102 420618 96134 421174
rect 95514 385174 96134 420618
rect 95514 384618 95546 385174
rect 96102 384618 96134 385174
rect 95514 349174 96134 384618
rect 95514 348618 95546 349174
rect 96102 348618 96134 349174
rect 95514 313174 96134 348618
rect 95514 312618 95546 313174
rect 96102 312618 96134 313174
rect 95514 277174 96134 312618
rect 95514 276618 95546 277174
rect 96102 276618 96134 277174
rect 95514 241174 96134 276618
rect 95514 240618 95546 241174
rect 96102 240618 96134 241174
rect 95514 205174 96134 240618
rect 95514 204618 95546 205174
rect 96102 204618 96134 205174
rect 95514 169174 96134 204618
rect 95514 168618 95546 169174
rect 96102 168618 96134 169174
rect 95514 133174 96134 168618
rect 95514 132618 95546 133174
rect 96102 132618 96134 133174
rect 95514 97174 96134 132618
rect 95514 96618 95546 97174
rect 96102 96618 96134 97174
rect 95514 61174 96134 96618
rect 95514 60618 95546 61174
rect 96102 60618 96134 61174
rect 95514 25174 96134 60618
rect 95514 24618 95546 25174
rect 96102 24618 96134 25174
rect 95514 -3226 96134 24618
rect 95514 -3782 95546 -3226
rect 96102 -3782 96134 -3226
rect 95514 -3814 96134 -3782
rect 99234 676894 99854 709082
rect 99234 676338 99266 676894
rect 99822 676338 99854 676894
rect 99234 640894 99854 676338
rect 99234 640338 99266 640894
rect 99822 640338 99854 640894
rect 99234 604894 99854 640338
rect 99234 604338 99266 604894
rect 99822 604338 99854 604894
rect 99234 568894 99854 604338
rect 99234 568338 99266 568894
rect 99822 568338 99854 568894
rect 99234 532894 99854 568338
rect 99234 532338 99266 532894
rect 99822 532338 99854 532894
rect 99234 496894 99854 532338
rect 99234 496338 99266 496894
rect 99822 496338 99854 496894
rect 99234 460894 99854 496338
rect 99234 460338 99266 460894
rect 99822 460338 99854 460894
rect 99234 424894 99854 460338
rect 99234 424338 99266 424894
rect 99822 424338 99854 424894
rect 99234 388894 99854 424338
rect 99234 388338 99266 388894
rect 99822 388338 99854 388894
rect 99234 352894 99854 388338
rect 99234 352338 99266 352894
rect 99822 352338 99854 352894
rect 99234 316894 99854 352338
rect 99234 316338 99266 316894
rect 99822 316338 99854 316894
rect 99234 280894 99854 316338
rect 99234 280338 99266 280894
rect 99822 280338 99854 280894
rect 99234 244894 99854 280338
rect 99234 244338 99266 244894
rect 99822 244338 99854 244894
rect 99234 208894 99854 244338
rect 99234 208338 99266 208894
rect 99822 208338 99854 208894
rect 99234 172894 99854 208338
rect 99234 172338 99266 172894
rect 99822 172338 99854 172894
rect 99234 136894 99854 172338
rect 99234 136338 99266 136894
rect 99822 136338 99854 136894
rect 99234 100894 99854 136338
rect 99234 100338 99266 100894
rect 99822 100338 99854 100894
rect 99234 64894 99854 100338
rect 99234 64338 99266 64894
rect 99822 64338 99854 64894
rect 99234 28894 99854 64338
rect 99234 28338 99266 28894
rect 99822 28338 99854 28894
rect 99234 -5146 99854 28338
rect 99234 -5702 99266 -5146
rect 99822 -5702 99854 -5146
rect 99234 -5734 99854 -5702
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710042 120986 710598
rect 121542 710042 121574 710598
rect 117234 708678 117854 709670
rect 117234 708122 117266 708678
rect 117822 708122 117854 708678
rect 113514 706758 114134 707750
rect 113514 706202 113546 706758
rect 114102 706202 114134 706758
rect 102954 680058 102986 680614
rect 103542 680058 103574 680614
rect 102954 644614 103574 680058
rect 102954 644058 102986 644614
rect 103542 644058 103574 644614
rect 102954 608614 103574 644058
rect 102954 608058 102986 608614
rect 103542 608058 103574 608614
rect 102954 572614 103574 608058
rect 102954 572058 102986 572614
rect 103542 572058 103574 572614
rect 102954 536614 103574 572058
rect 102954 536058 102986 536614
rect 103542 536058 103574 536614
rect 102954 500614 103574 536058
rect 102954 500058 102986 500614
rect 103542 500058 103574 500614
rect 102954 464614 103574 500058
rect 102954 464058 102986 464614
rect 103542 464058 103574 464614
rect 102954 428614 103574 464058
rect 102954 428058 102986 428614
rect 103542 428058 103574 428614
rect 102954 392614 103574 428058
rect 102954 392058 102986 392614
rect 103542 392058 103574 392614
rect 102954 356614 103574 392058
rect 102954 356058 102986 356614
rect 103542 356058 103574 356614
rect 102954 320614 103574 356058
rect 102954 320058 102986 320614
rect 103542 320058 103574 320614
rect 102954 284614 103574 320058
rect 102954 284058 102986 284614
rect 103542 284058 103574 284614
rect 102954 248614 103574 284058
rect 102954 248058 102986 248614
rect 103542 248058 103574 248614
rect 102954 212614 103574 248058
rect 102954 212058 102986 212614
rect 103542 212058 103574 212614
rect 102954 176614 103574 212058
rect 102954 176058 102986 176614
rect 103542 176058 103574 176614
rect 102954 140614 103574 176058
rect 102954 140058 102986 140614
rect 103542 140058 103574 140614
rect 102954 104614 103574 140058
rect 102954 104058 102986 104614
rect 103542 104058 103574 104614
rect 102954 68614 103574 104058
rect 102954 68058 102986 68614
rect 103542 68058 103574 68614
rect 102954 32614 103574 68058
rect 102954 32058 102986 32614
rect 103542 32058 103574 32614
rect 84954 -6662 84986 -6106
rect 85542 -6662 85574 -6106
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 704838 110414 705830
rect 109794 704282 109826 704838
rect 110382 704282 110414 704838
rect 109794 687454 110414 704282
rect 109794 686898 109826 687454
rect 110382 686898 110414 687454
rect 109794 651454 110414 686898
rect 109794 650898 109826 651454
rect 110382 650898 110414 651454
rect 109794 615454 110414 650898
rect 109794 614898 109826 615454
rect 110382 614898 110414 615454
rect 109794 579454 110414 614898
rect 109794 578898 109826 579454
rect 110382 578898 110414 579454
rect 109794 543454 110414 578898
rect 109794 542898 109826 543454
rect 110382 542898 110414 543454
rect 109794 507454 110414 542898
rect 109794 506898 109826 507454
rect 110382 506898 110414 507454
rect 109794 471454 110414 506898
rect 109794 470898 109826 471454
rect 110382 470898 110414 471454
rect 109794 435454 110414 470898
rect 109794 434898 109826 435454
rect 110382 434898 110414 435454
rect 109794 399454 110414 434898
rect 109794 398898 109826 399454
rect 110382 398898 110414 399454
rect 109794 363454 110414 398898
rect 109794 362898 109826 363454
rect 110382 362898 110414 363454
rect 109794 327454 110414 362898
rect 109794 326898 109826 327454
rect 110382 326898 110414 327454
rect 109794 291454 110414 326898
rect 109794 290898 109826 291454
rect 110382 290898 110414 291454
rect 109794 255454 110414 290898
rect 109794 254898 109826 255454
rect 110382 254898 110414 255454
rect 109794 219454 110414 254898
rect 109794 218898 109826 219454
rect 110382 218898 110414 219454
rect 109794 183454 110414 218898
rect 109794 182898 109826 183454
rect 110382 182898 110414 183454
rect 109794 147454 110414 182898
rect 109794 146898 109826 147454
rect 110382 146898 110414 147454
rect 109794 111454 110414 146898
rect 109794 110898 109826 111454
rect 110382 110898 110414 111454
rect 109794 75454 110414 110898
rect 109794 74898 109826 75454
rect 110382 74898 110414 75454
rect 109794 39454 110414 74898
rect 109794 38898 109826 39454
rect 110382 38898 110414 39454
rect 109794 3454 110414 38898
rect 109794 2898 109826 3454
rect 110382 2898 110414 3454
rect 109794 -346 110414 2898
rect 109794 -902 109826 -346
rect 110382 -902 110414 -346
rect 109794 -1894 110414 -902
rect 113514 691174 114134 706202
rect 113514 690618 113546 691174
rect 114102 690618 114134 691174
rect 113514 655174 114134 690618
rect 113514 654618 113546 655174
rect 114102 654618 114134 655174
rect 113514 619174 114134 654618
rect 113514 618618 113546 619174
rect 114102 618618 114134 619174
rect 113514 583174 114134 618618
rect 113514 582618 113546 583174
rect 114102 582618 114134 583174
rect 113514 547174 114134 582618
rect 113514 546618 113546 547174
rect 114102 546618 114134 547174
rect 113514 511174 114134 546618
rect 113514 510618 113546 511174
rect 114102 510618 114134 511174
rect 113514 475174 114134 510618
rect 113514 474618 113546 475174
rect 114102 474618 114134 475174
rect 113514 439174 114134 474618
rect 113514 438618 113546 439174
rect 114102 438618 114134 439174
rect 113514 403174 114134 438618
rect 113514 402618 113546 403174
rect 114102 402618 114134 403174
rect 113514 367174 114134 402618
rect 113514 366618 113546 367174
rect 114102 366618 114134 367174
rect 113514 331174 114134 366618
rect 113514 330618 113546 331174
rect 114102 330618 114134 331174
rect 113514 295174 114134 330618
rect 113514 294618 113546 295174
rect 114102 294618 114134 295174
rect 113514 259174 114134 294618
rect 113514 258618 113546 259174
rect 114102 258618 114134 259174
rect 113514 223174 114134 258618
rect 113514 222618 113546 223174
rect 114102 222618 114134 223174
rect 113514 187174 114134 222618
rect 113514 186618 113546 187174
rect 114102 186618 114134 187174
rect 113514 151174 114134 186618
rect 113514 150618 113546 151174
rect 114102 150618 114134 151174
rect 113514 115174 114134 150618
rect 113514 114618 113546 115174
rect 114102 114618 114134 115174
rect 113514 79174 114134 114618
rect 113514 78618 113546 79174
rect 114102 78618 114134 79174
rect 113514 43174 114134 78618
rect 113514 42618 113546 43174
rect 114102 42618 114134 43174
rect 113514 7174 114134 42618
rect 113514 6618 113546 7174
rect 114102 6618 114134 7174
rect 113514 -2266 114134 6618
rect 113514 -2822 113546 -2266
rect 114102 -2822 114134 -2266
rect 113514 -3814 114134 -2822
rect 117234 694894 117854 708122
rect 117234 694338 117266 694894
rect 117822 694338 117854 694894
rect 117234 658894 117854 694338
rect 117234 658338 117266 658894
rect 117822 658338 117854 658894
rect 117234 622894 117854 658338
rect 117234 622338 117266 622894
rect 117822 622338 117854 622894
rect 117234 586894 117854 622338
rect 117234 586338 117266 586894
rect 117822 586338 117854 586894
rect 117234 550894 117854 586338
rect 117234 550338 117266 550894
rect 117822 550338 117854 550894
rect 117234 514894 117854 550338
rect 117234 514338 117266 514894
rect 117822 514338 117854 514894
rect 117234 478894 117854 514338
rect 117234 478338 117266 478894
rect 117822 478338 117854 478894
rect 117234 442894 117854 478338
rect 117234 442338 117266 442894
rect 117822 442338 117854 442894
rect 117234 406894 117854 442338
rect 117234 406338 117266 406894
rect 117822 406338 117854 406894
rect 117234 370894 117854 406338
rect 117234 370338 117266 370894
rect 117822 370338 117854 370894
rect 117234 334894 117854 370338
rect 117234 334338 117266 334894
rect 117822 334338 117854 334894
rect 117234 298894 117854 334338
rect 117234 298338 117266 298894
rect 117822 298338 117854 298894
rect 117234 262894 117854 298338
rect 117234 262338 117266 262894
rect 117822 262338 117854 262894
rect 117234 226894 117854 262338
rect 117234 226338 117266 226894
rect 117822 226338 117854 226894
rect 117234 190894 117854 226338
rect 117234 190338 117266 190894
rect 117822 190338 117854 190894
rect 117234 154894 117854 190338
rect 117234 154338 117266 154894
rect 117822 154338 117854 154894
rect 117234 118894 117854 154338
rect 117234 118338 117266 118894
rect 117822 118338 117854 118894
rect 117234 82894 117854 118338
rect 117234 82338 117266 82894
rect 117822 82338 117854 82894
rect 117234 46894 117854 82338
rect 117234 46338 117266 46894
rect 117822 46338 117854 46894
rect 117234 10894 117854 46338
rect 117234 10338 117266 10894
rect 117822 10338 117854 10894
rect 117234 -4186 117854 10338
rect 117234 -4742 117266 -4186
rect 117822 -4742 117854 -4186
rect 117234 -5734 117854 -4742
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711002 138986 711558
rect 139542 711002 139574 711558
rect 135234 709638 135854 709670
rect 135234 709082 135266 709638
rect 135822 709082 135854 709638
rect 131514 707718 132134 707750
rect 131514 707162 131546 707718
rect 132102 707162 132134 707718
rect 120954 698058 120986 698614
rect 121542 698058 121574 698614
rect 120954 662614 121574 698058
rect 120954 662058 120986 662614
rect 121542 662058 121574 662614
rect 120954 626614 121574 662058
rect 120954 626058 120986 626614
rect 121542 626058 121574 626614
rect 120954 590614 121574 626058
rect 120954 590058 120986 590614
rect 121542 590058 121574 590614
rect 120954 554614 121574 590058
rect 120954 554058 120986 554614
rect 121542 554058 121574 554614
rect 120954 518614 121574 554058
rect 120954 518058 120986 518614
rect 121542 518058 121574 518614
rect 120954 482614 121574 518058
rect 120954 482058 120986 482614
rect 121542 482058 121574 482614
rect 120954 446614 121574 482058
rect 120954 446058 120986 446614
rect 121542 446058 121574 446614
rect 120954 410614 121574 446058
rect 120954 410058 120986 410614
rect 121542 410058 121574 410614
rect 120954 374614 121574 410058
rect 120954 374058 120986 374614
rect 121542 374058 121574 374614
rect 120954 338614 121574 374058
rect 120954 338058 120986 338614
rect 121542 338058 121574 338614
rect 120954 302614 121574 338058
rect 120954 302058 120986 302614
rect 121542 302058 121574 302614
rect 120954 266614 121574 302058
rect 120954 266058 120986 266614
rect 121542 266058 121574 266614
rect 120954 230614 121574 266058
rect 120954 230058 120986 230614
rect 121542 230058 121574 230614
rect 120954 194614 121574 230058
rect 120954 194058 120986 194614
rect 121542 194058 121574 194614
rect 120954 158614 121574 194058
rect 120954 158058 120986 158614
rect 121542 158058 121574 158614
rect 120954 122614 121574 158058
rect 120954 122058 120986 122614
rect 121542 122058 121574 122614
rect 120954 86614 121574 122058
rect 120954 86058 120986 86614
rect 121542 86058 121574 86614
rect 120954 50614 121574 86058
rect 120954 50058 120986 50614
rect 121542 50058 121574 50614
rect 120954 14614 121574 50058
rect 120954 14058 120986 14614
rect 121542 14058 121574 14614
rect 102954 -7622 102986 -7066
rect 103542 -7622 103574 -7066
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 705798 128414 705830
rect 127794 705242 127826 705798
rect 128382 705242 128414 705798
rect 127794 669454 128414 705242
rect 127794 668898 127826 669454
rect 128382 668898 128414 669454
rect 127794 633454 128414 668898
rect 127794 632898 127826 633454
rect 128382 632898 128414 633454
rect 127794 597454 128414 632898
rect 127794 596898 127826 597454
rect 128382 596898 128414 597454
rect 127794 561454 128414 596898
rect 127794 560898 127826 561454
rect 128382 560898 128414 561454
rect 127794 525454 128414 560898
rect 127794 524898 127826 525454
rect 128382 524898 128414 525454
rect 127794 489454 128414 524898
rect 127794 488898 127826 489454
rect 128382 488898 128414 489454
rect 127794 453454 128414 488898
rect 127794 452898 127826 453454
rect 128382 452898 128414 453454
rect 127794 417454 128414 452898
rect 127794 416898 127826 417454
rect 128382 416898 128414 417454
rect 127794 381454 128414 416898
rect 127794 380898 127826 381454
rect 128382 380898 128414 381454
rect 127794 345454 128414 380898
rect 127794 344898 127826 345454
rect 128382 344898 128414 345454
rect 127794 309454 128414 344898
rect 127794 308898 127826 309454
rect 128382 308898 128414 309454
rect 127794 273454 128414 308898
rect 127794 272898 127826 273454
rect 128382 272898 128414 273454
rect 127794 237454 128414 272898
rect 127794 236898 127826 237454
rect 128382 236898 128414 237454
rect 127794 201454 128414 236898
rect 127794 200898 127826 201454
rect 128382 200898 128414 201454
rect 127794 165454 128414 200898
rect 127794 164898 127826 165454
rect 128382 164898 128414 165454
rect 127794 129454 128414 164898
rect 127794 128898 127826 129454
rect 128382 128898 128414 129454
rect 127794 93454 128414 128898
rect 127794 92898 127826 93454
rect 128382 92898 128414 93454
rect 127794 57454 128414 92898
rect 127794 56898 127826 57454
rect 128382 56898 128414 57454
rect 127794 21454 128414 56898
rect 127794 20898 127826 21454
rect 128382 20898 128414 21454
rect 127794 -1306 128414 20898
rect 127794 -1862 127826 -1306
rect 128382 -1862 128414 -1306
rect 127794 -1894 128414 -1862
rect 131514 673174 132134 707162
rect 131514 672618 131546 673174
rect 132102 672618 132134 673174
rect 131514 637174 132134 672618
rect 131514 636618 131546 637174
rect 132102 636618 132134 637174
rect 131514 601174 132134 636618
rect 131514 600618 131546 601174
rect 132102 600618 132134 601174
rect 131514 565174 132134 600618
rect 131514 564618 131546 565174
rect 132102 564618 132134 565174
rect 131514 529174 132134 564618
rect 131514 528618 131546 529174
rect 132102 528618 132134 529174
rect 131514 493174 132134 528618
rect 131514 492618 131546 493174
rect 132102 492618 132134 493174
rect 131514 457174 132134 492618
rect 131514 456618 131546 457174
rect 132102 456618 132134 457174
rect 131514 421174 132134 456618
rect 131514 420618 131546 421174
rect 132102 420618 132134 421174
rect 131514 385174 132134 420618
rect 131514 384618 131546 385174
rect 132102 384618 132134 385174
rect 131514 349174 132134 384618
rect 131514 348618 131546 349174
rect 132102 348618 132134 349174
rect 131514 313174 132134 348618
rect 131514 312618 131546 313174
rect 132102 312618 132134 313174
rect 131514 277174 132134 312618
rect 131514 276618 131546 277174
rect 132102 276618 132134 277174
rect 131514 241174 132134 276618
rect 131514 240618 131546 241174
rect 132102 240618 132134 241174
rect 131514 205174 132134 240618
rect 131514 204618 131546 205174
rect 132102 204618 132134 205174
rect 131514 169174 132134 204618
rect 131514 168618 131546 169174
rect 132102 168618 132134 169174
rect 131514 133174 132134 168618
rect 131514 132618 131546 133174
rect 132102 132618 132134 133174
rect 131514 97174 132134 132618
rect 131514 96618 131546 97174
rect 132102 96618 132134 97174
rect 131514 61174 132134 96618
rect 131514 60618 131546 61174
rect 132102 60618 132134 61174
rect 131514 25174 132134 60618
rect 131514 24618 131546 25174
rect 132102 24618 132134 25174
rect 131514 -3226 132134 24618
rect 131514 -3782 131546 -3226
rect 132102 -3782 132134 -3226
rect 131514 -3814 132134 -3782
rect 135234 676894 135854 709082
rect 135234 676338 135266 676894
rect 135822 676338 135854 676894
rect 135234 640894 135854 676338
rect 135234 640338 135266 640894
rect 135822 640338 135854 640894
rect 135234 604894 135854 640338
rect 135234 604338 135266 604894
rect 135822 604338 135854 604894
rect 135234 568894 135854 604338
rect 135234 568338 135266 568894
rect 135822 568338 135854 568894
rect 135234 532894 135854 568338
rect 135234 532338 135266 532894
rect 135822 532338 135854 532894
rect 135234 496894 135854 532338
rect 135234 496338 135266 496894
rect 135822 496338 135854 496894
rect 135234 460894 135854 496338
rect 135234 460338 135266 460894
rect 135822 460338 135854 460894
rect 135234 424894 135854 460338
rect 135234 424338 135266 424894
rect 135822 424338 135854 424894
rect 135234 388894 135854 424338
rect 135234 388338 135266 388894
rect 135822 388338 135854 388894
rect 135234 352894 135854 388338
rect 135234 352338 135266 352894
rect 135822 352338 135854 352894
rect 135234 316894 135854 352338
rect 135234 316338 135266 316894
rect 135822 316338 135854 316894
rect 135234 280894 135854 316338
rect 135234 280338 135266 280894
rect 135822 280338 135854 280894
rect 135234 244894 135854 280338
rect 135234 244338 135266 244894
rect 135822 244338 135854 244894
rect 135234 208894 135854 244338
rect 135234 208338 135266 208894
rect 135822 208338 135854 208894
rect 135234 172894 135854 208338
rect 135234 172338 135266 172894
rect 135822 172338 135854 172894
rect 135234 136894 135854 172338
rect 135234 136338 135266 136894
rect 135822 136338 135854 136894
rect 135234 100894 135854 136338
rect 135234 100338 135266 100894
rect 135822 100338 135854 100894
rect 135234 64894 135854 100338
rect 135234 64338 135266 64894
rect 135822 64338 135854 64894
rect 135234 28894 135854 64338
rect 135234 28338 135266 28894
rect 135822 28338 135854 28894
rect 135234 -5146 135854 28338
rect 135234 -5702 135266 -5146
rect 135822 -5702 135854 -5146
rect 135234 -5734 135854 -5702
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710042 156986 710598
rect 157542 710042 157574 710598
rect 153234 708678 153854 709670
rect 153234 708122 153266 708678
rect 153822 708122 153854 708678
rect 149514 706758 150134 707750
rect 149514 706202 149546 706758
rect 150102 706202 150134 706758
rect 138954 680058 138986 680614
rect 139542 680058 139574 680614
rect 138954 644614 139574 680058
rect 138954 644058 138986 644614
rect 139542 644058 139574 644614
rect 138954 608614 139574 644058
rect 138954 608058 138986 608614
rect 139542 608058 139574 608614
rect 138954 572614 139574 608058
rect 138954 572058 138986 572614
rect 139542 572058 139574 572614
rect 138954 536614 139574 572058
rect 138954 536058 138986 536614
rect 139542 536058 139574 536614
rect 138954 500614 139574 536058
rect 138954 500058 138986 500614
rect 139542 500058 139574 500614
rect 138954 464614 139574 500058
rect 138954 464058 138986 464614
rect 139542 464058 139574 464614
rect 138954 428614 139574 464058
rect 138954 428058 138986 428614
rect 139542 428058 139574 428614
rect 138954 392614 139574 428058
rect 138954 392058 138986 392614
rect 139542 392058 139574 392614
rect 138954 356614 139574 392058
rect 138954 356058 138986 356614
rect 139542 356058 139574 356614
rect 138954 320614 139574 356058
rect 138954 320058 138986 320614
rect 139542 320058 139574 320614
rect 138954 284614 139574 320058
rect 138954 284058 138986 284614
rect 139542 284058 139574 284614
rect 138954 248614 139574 284058
rect 138954 248058 138986 248614
rect 139542 248058 139574 248614
rect 138954 212614 139574 248058
rect 138954 212058 138986 212614
rect 139542 212058 139574 212614
rect 138954 176614 139574 212058
rect 138954 176058 138986 176614
rect 139542 176058 139574 176614
rect 138954 140614 139574 176058
rect 138954 140058 138986 140614
rect 139542 140058 139574 140614
rect 138954 104614 139574 140058
rect 138954 104058 138986 104614
rect 139542 104058 139574 104614
rect 138954 68614 139574 104058
rect 138954 68058 138986 68614
rect 139542 68058 139574 68614
rect 138954 32614 139574 68058
rect 138954 32058 138986 32614
rect 139542 32058 139574 32614
rect 120954 -6662 120986 -6106
rect 121542 -6662 121574 -6106
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 704838 146414 705830
rect 145794 704282 145826 704838
rect 146382 704282 146414 704838
rect 145794 687454 146414 704282
rect 145794 686898 145826 687454
rect 146382 686898 146414 687454
rect 145794 651454 146414 686898
rect 145794 650898 145826 651454
rect 146382 650898 146414 651454
rect 145794 615454 146414 650898
rect 145794 614898 145826 615454
rect 146382 614898 146414 615454
rect 145794 579454 146414 614898
rect 145794 578898 145826 579454
rect 146382 578898 146414 579454
rect 145794 543454 146414 578898
rect 145794 542898 145826 543454
rect 146382 542898 146414 543454
rect 145794 507454 146414 542898
rect 145794 506898 145826 507454
rect 146382 506898 146414 507454
rect 145794 471454 146414 506898
rect 145794 470898 145826 471454
rect 146382 470898 146414 471454
rect 145794 435454 146414 470898
rect 145794 434898 145826 435454
rect 146382 434898 146414 435454
rect 145794 399454 146414 434898
rect 145794 398898 145826 399454
rect 146382 398898 146414 399454
rect 145794 363454 146414 398898
rect 145794 362898 145826 363454
rect 146382 362898 146414 363454
rect 145794 327454 146414 362898
rect 145794 326898 145826 327454
rect 146382 326898 146414 327454
rect 145794 291454 146414 326898
rect 145794 290898 145826 291454
rect 146382 290898 146414 291454
rect 145794 255454 146414 290898
rect 145794 254898 145826 255454
rect 146382 254898 146414 255454
rect 145794 219454 146414 254898
rect 145794 218898 145826 219454
rect 146382 218898 146414 219454
rect 145794 183454 146414 218898
rect 145794 182898 145826 183454
rect 146382 182898 146414 183454
rect 145794 147454 146414 182898
rect 145794 146898 145826 147454
rect 146382 146898 146414 147454
rect 145794 111454 146414 146898
rect 145794 110898 145826 111454
rect 146382 110898 146414 111454
rect 145794 75454 146414 110898
rect 145794 74898 145826 75454
rect 146382 74898 146414 75454
rect 145794 39454 146414 74898
rect 145794 38898 145826 39454
rect 146382 38898 146414 39454
rect 145794 3454 146414 38898
rect 145794 2898 145826 3454
rect 146382 2898 146414 3454
rect 145794 -346 146414 2898
rect 145794 -902 145826 -346
rect 146382 -902 146414 -346
rect 145794 -1894 146414 -902
rect 149514 691174 150134 706202
rect 149514 690618 149546 691174
rect 150102 690618 150134 691174
rect 149514 655174 150134 690618
rect 149514 654618 149546 655174
rect 150102 654618 150134 655174
rect 149514 619174 150134 654618
rect 149514 618618 149546 619174
rect 150102 618618 150134 619174
rect 149514 583174 150134 618618
rect 149514 582618 149546 583174
rect 150102 582618 150134 583174
rect 149514 547174 150134 582618
rect 149514 546618 149546 547174
rect 150102 546618 150134 547174
rect 149514 511174 150134 546618
rect 149514 510618 149546 511174
rect 150102 510618 150134 511174
rect 149514 475174 150134 510618
rect 149514 474618 149546 475174
rect 150102 474618 150134 475174
rect 149514 439174 150134 474618
rect 149514 438618 149546 439174
rect 150102 438618 150134 439174
rect 149514 403174 150134 438618
rect 149514 402618 149546 403174
rect 150102 402618 150134 403174
rect 149514 367174 150134 402618
rect 149514 366618 149546 367174
rect 150102 366618 150134 367174
rect 149514 331174 150134 366618
rect 149514 330618 149546 331174
rect 150102 330618 150134 331174
rect 149514 295174 150134 330618
rect 149514 294618 149546 295174
rect 150102 294618 150134 295174
rect 149514 259174 150134 294618
rect 149514 258618 149546 259174
rect 150102 258618 150134 259174
rect 149514 223174 150134 258618
rect 149514 222618 149546 223174
rect 150102 222618 150134 223174
rect 149514 187174 150134 222618
rect 149514 186618 149546 187174
rect 150102 186618 150134 187174
rect 149514 151174 150134 186618
rect 149514 150618 149546 151174
rect 150102 150618 150134 151174
rect 149514 115174 150134 150618
rect 149514 114618 149546 115174
rect 150102 114618 150134 115174
rect 149514 79174 150134 114618
rect 149514 78618 149546 79174
rect 150102 78618 150134 79174
rect 149514 43174 150134 78618
rect 149514 42618 149546 43174
rect 150102 42618 150134 43174
rect 149514 7174 150134 42618
rect 149514 6618 149546 7174
rect 150102 6618 150134 7174
rect 149514 -2266 150134 6618
rect 149514 -2822 149546 -2266
rect 150102 -2822 150134 -2266
rect 149514 -3814 150134 -2822
rect 153234 694894 153854 708122
rect 153234 694338 153266 694894
rect 153822 694338 153854 694894
rect 153234 658894 153854 694338
rect 153234 658338 153266 658894
rect 153822 658338 153854 658894
rect 153234 622894 153854 658338
rect 153234 622338 153266 622894
rect 153822 622338 153854 622894
rect 153234 586894 153854 622338
rect 153234 586338 153266 586894
rect 153822 586338 153854 586894
rect 153234 550894 153854 586338
rect 153234 550338 153266 550894
rect 153822 550338 153854 550894
rect 153234 514894 153854 550338
rect 153234 514338 153266 514894
rect 153822 514338 153854 514894
rect 153234 478894 153854 514338
rect 153234 478338 153266 478894
rect 153822 478338 153854 478894
rect 153234 442894 153854 478338
rect 153234 442338 153266 442894
rect 153822 442338 153854 442894
rect 153234 406894 153854 442338
rect 153234 406338 153266 406894
rect 153822 406338 153854 406894
rect 153234 370894 153854 406338
rect 153234 370338 153266 370894
rect 153822 370338 153854 370894
rect 153234 334894 153854 370338
rect 153234 334338 153266 334894
rect 153822 334338 153854 334894
rect 153234 298894 153854 334338
rect 153234 298338 153266 298894
rect 153822 298338 153854 298894
rect 153234 262894 153854 298338
rect 153234 262338 153266 262894
rect 153822 262338 153854 262894
rect 153234 226894 153854 262338
rect 153234 226338 153266 226894
rect 153822 226338 153854 226894
rect 153234 190894 153854 226338
rect 153234 190338 153266 190894
rect 153822 190338 153854 190894
rect 153234 154894 153854 190338
rect 153234 154338 153266 154894
rect 153822 154338 153854 154894
rect 153234 118894 153854 154338
rect 153234 118338 153266 118894
rect 153822 118338 153854 118894
rect 153234 82894 153854 118338
rect 153234 82338 153266 82894
rect 153822 82338 153854 82894
rect 153234 46894 153854 82338
rect 153234 46338 153266 46894
rect 153822 46338 153854 46894
rect 153234 10894 153854 46338
rect 153234 10338 153266 10894
rect 153822 10338 153854 10894
rect 153234 -4186 153854 10338
rect 153234 -4742 153266 -4186
rect 153822 -4742 153854 -4186
rect 153234 -5734 153854 -4742
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711002 174986 711558
rect 175542 711002 175574 711558
rect 171234 709638 171854 709670
rect 171234 709082 171266 709638
rect 171822 709082 171854 709638
rect 167514 707718 168134 707750
rect 167514 707162 167546 707718
rect 168102 707162 168134 707718
rect 156954 698058 156986 698614
rect 157542 698058 157574 698614
rect 156954 662614 157574 698058
rect 156954 662058 156986 662614
rect 157542 662058 157574 662614
rect 156954 626614 157574 662058
rect 156954 626058 156986 626614
rect 157542 626058 157574 626614
rect 156954 590614 157574 626058
rect 156954 590058 156986 590614
rect 157542 590058 157574 590614
rect 156954 554614 157574 590058
rect 156954 554058 156986 554614
rect 157542 554058 157574 554614
rect 156954 518614 157574 554058
rect 156954 518058 156986 518614
rect 157542 518058 157574 518614
rect 156954 482614 157574 518058
rect 156954 482058 156986 482614
rect 157542 482058 157574 482614
rect 156954 446614 157574 482058
rect 156954 446058 156986 446614
rect 157542 446058 157574 446614
rect 156954 410614 157574 446058
rect 156954 410058 156986 410614
rect 157542 410058 157574 410614
rect 156954 374614 157574 410058
rect 156954 374058 156986 374614
rect 157542 374058 157574 374614
rect 156954 338614 157574 374058
rect 156954 338058 156986 338614
rect 157542 338058 157574 338614
rect 156954 302614 157574 338058
rect 156954 302058 156986 302614
rect 157542 302058 157574 302614
rect 156954 266614 157574 302058
rect 156954 266058 156986 266614
rect 157542 266058 157574 266614
rect 156954 230614 157574 266058
rect 156954 230058 156986 230614
rect 157542 230058 157574 230614
rect 156954 194614 157574 230058
rect 156954 194058 156986 194614
rect 157542 194058 157574 194614
rect 156954 158614 157574 194058
rect 156954 158058 156986 158614
rect 157542 158058 157574 158614
rect 156954 122614 157574 158058
rect 156954 122058 156986 122614
rect 157542 122058 157574 122614
rect 156954 86614 157574 122058
rect 156954 86058 156986 86614
rect 157542 86058 157574 86614
rect 156954 50614 157574 86058
rect 156954 50058 156986 50614
rect 157542 50058 157574 50614
rect 156954 14614 157574 50058
rect 156954 14058 156986 14614
rect 157542 14058 157574 14614
rect 138954 -7622 138986 -7066
rect 139542 -7622 139574 -7066
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 705798 164414 705830
rect 163794 705242 163826 705798
rect 164382 705242 164414 705798
rect 163794 669454 164414 705242
rect 163794 668898 163826 669454
rect 164382 668898 164414 669454
rect 163794 633454 164414 668898
rect 163794 632898 163826 633454
rect 164382 632898 164414 633454
rect 163794 597454 164414 632898
rect 163794 596898 163826 597454
rect 164382 596898 164414 597454
rect 163794 561454 164414 596898
rect 163794 560898 163826 561454
rect 164382 560898 164414 561454
rect 163794 525454 164414 560898
rect 163794 524898 163826 525454
rect 164382 524898 164414 525454
rect 163794 489454 164414 524898
rect 163794 488898 163826 489454
rect 164382 488898 164414 489454
rect 163794 453454 164414 488898
rect 163794 452898 163826 453454
rect 164382 452898 164414 453454
rect 163794 417454 164414 452898
rect 163794 416898 163826 417454
rect 164382 416898 164414 417454
rect 163794 381454 164414 416898
rect 163794 380898 163826 381454
rect 164382 380898 164414 381454
rect 163794 345454 164414 380898
rect 163794 344898 163826 345454
rect 164382 344898 164414 345454
rect 163794 309454 164414 344898
rect 163794 308898 163826 309454
rect 164382 308898 164414 309454
rect 163794 273454 164414 308898
rect 163794 272898 163826 273454
rect 164382 272898 164414 273454
rect 163794 237454 164414 272898
rect 163794 236898 163826 237454
rect 164382 236898 164414 237454
rect 163794 201454 164414 236898
rect 163794 200898 163826 201454
rect 164382 200898 164414 201454
rect 163794 165454 164414 200898
rect 163794 164898 163826 165454
rect 164382 164898 164414 165454
rect 163794 129454 164414 164898
rect 163794 128898 163826 129454
rect 164382 128898 164414 129454
rect 163794 93454 164414 128898
rect 163794 92898 163826 93454
rect 164382 92898 164414 93454
rect 163794 57454 164414 92898
rect 163794 56898 163826 57454
rect 164382 56898 164414 57454
rect 163794 21454 164414 56898
rect 163794 20898 163826 21454
rect 164382 20898 164414 21454
rect 163794 -1306 164414 20898
rect 163794 -1862 163826 -1306
rect 164382 -1862 164414 -1306
rect 163794 -1894 164414 -1862
rect 167514 673174 168134 707162
rect 167514 672618 167546 673174
rect 168102 672618 168134 673174
rect 167514 637174 168134 672618
rect 167514 636618 167546 637174
rect 168102 636618 168134 637174
rect 167514 601174 168134 636618
rect 167514 600618 167546 601174
rect 168102 600618 168134 601174
rect 167514 565174 168134 600618
rect 167514 564618 167546 565174
rect 168102 564618 168134 565174
rect 167514 529174 168134 564618
rect 167514 528618 167546 529174
rect 168102 528618 168134 529174
rect 167514 493174 168134 528618
rect 167514 492618 167546 493174
rect 168102 492618 168134 493174
rect 167514 457174 168134 492618
rect 167514 456618 167546 457174
rect 168102 456618 168134 457174
rect 167514 421174 168134 456618
rect 167514 420618 167546 421174
rect 168102 420618 168134 421174
rect 167514 385174 168134 420618
rect 167514 384618 167546 385174
rect 168102 384618 168134 385174
rect 167514 349174 168134 384618
rect 167514 348618 167546 349174
rect 168102 348618 168134 349174
rect 167514 313174 168134 348618
rect 167514 312618 167546 313174
rect 168102 312618 168134 313174
rect 167514 277174 168134 312618
rect 167514 276618 167546 277174
rect 168102 276618 168134 277174
rect 167514 241174 168134 276618
rect 167514 240618 167546 241174
rect 168102 240618 168134 241174
rect 167514 205174 168134 240618
rect 167514 204618 167546 205174
rect 168102 204618 168134 205174
rect 167514 169174 168134 204618
rect 167514 168618 167546 169174
rect 168102 168618 168134 169174
rect 167514 133174 168134 168618
rect 167514 132618 167546 133174
rect 168102 132618 168134 133174
rect 167514 97174 168134 132618
rect 167514 96618 167546 97174
rect 168102 96618 168134 97174
rect 167514 61174 168134 96618
rect 167514 60618 167546 61174
rect 168102 60618 168134 61174
rect 167514 25174 168134 60618
rect 167514 24618 167546 25174
rect 168102 24618 168134 25174
rect 167514 -3226 168134 24618
rect 167514 -3782 167546 -3226
rect 168102 -3782 168134 -3226
rect 167514 -3814 168134 -3782
rect 171234 676894 171854 709082
rect 171234 676338 171266 676894
rect 171822 676338 171854 676894
rect 171234 640894 171854 676338
rect 171234 640338 171266 640894
rect 171822 640338 171854 640894
rect 171234 604894 171854 640338
rect 171234 604338 171266 604894
rect 171822 604338 171854 604894
rect 171234 568894 171854 604338
rect 171234 568338 171266 568894
rect 171822 568338 171854 568894
rect 171234 532894 171854 568338
rect 171234 532338 171266 532894
rect 171822 532338 171854 532894
rect 171234 496894 171854 532338
rect 171234 496338 171266 496894
rect 171822 496338 171854 496894
rect 171234 460894 171854 496338
rect 171234 460338 171266 460894
rect 171822 460338 171854 460894
rect 171234 424894 171854 460338
rect 171234 424338 171266 424894
rect 171822 424338 171854 424894
rect 171234 388894 171854 424338
rect 171234 388338 171266 388894
rect 171822 388338 171854 388894
rect 171234 352894 171854 388338
rect 171234 352338 171266 352894
rect 171822 352338 171854 352894
rect 171234 316894 171854 352338
rect 171234 316338 171266 316894
rect 171822 316338 171854 316894
rect 171234 280894 171854 316338
rect 171234 280338 171266 280894
rect 171822 280338 171854 280894
rect 171234 244894 171854 280338
rect 171234 244338 171266 244894
rect 171822 244338 171854 244894
rect 171234 208894 171854 244338
rect 171234 208338 171266 208894
rect 171822 208338 171854 208894
rect 171234 172894 171854 208338
rect 171234 172338 171266 172894
rect 171822 172338 171854 172894
rect 171234 136894 171854 172338
rect 171234 136338 171266 136894
rect 171822 136338 171854 136894
rect 171234 100894 171854 136338
rect 171234 100338 171266 100894
rect 171822 100338 171854 100894
rect 171234 64894 171854 100338
rect 171234 64338 171266 64894
rect 171822 64338 171854 64894
rect 171234 28894 171854 64338
rect 171234 28338 171266 28894
rect 171822 28338 171854 28894
rect 171234 -5146 171854 28338
rect 171234 -5702 171266 -5146
rect 171822 -5702 171854 -5146
rect 171234 -5734 171854 -5702
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710042 192986 710598
rect 193542 710042 193574 710598
rect 189234 708678 189854 709670
rect 189234 708122 189266 708678
rect 189822 708122 189854 708678
rect 185514 706758 186134 707750
rect 185514 706202 185546 706758
rect 186102 706202 186134 706758
rect 174954 680058 174986 680614
rect 175542 680058 175574 680614
rect 174954 644614 175574 680058
rect 174954 644058 174986 644614
rect 175542 644058 175574 644614
rect 174954 608614 175574 644058
rect 174954 608058 174986 608614
rect 175542 608058 175574 608614
rect 174954 572614 175574 608058
rect 174954 572058 174986 572614
rect 175542 572058 175574 572614
rect 174954 536614 175574 572058
rect 174954 536058 174986 536614
rect 175542 536058 175574 536614
rect 174954 500614 175574 536058
rect 174954 500058 174986 500614
rect 175542 500058 175574 500614
rect 174954 464614 175574 500058
rect 174954 464058 174986 464614
rect 175542 464058 175574 464614
rect 174954 428614 175574 464058
rect 174954 428058 174986 428614
rect 175542 428058 175574 428614
rect 174954 392614 175574 428058
rect 174954 392058 174986 392614
rect 175542 392058 175574 392614
rect 174954 356614 175574 392058
rect 174954 356058 174986 356614
rect 175542 356058 175574 356614
rect 174954 320614 175574 356058
rect 174954 320058 174986 320614
rect 175542 320058 175574 320614
rect 174954 284614 175574 320058
rect 174954 284058 174986 284614
rect 175542 284058 175574 284614
rect 174954 248614 175574 284058
rect 174954 248058 174986 248614
rect 175542 248058 175574 248614
rect 174954 212614 175574 248058
rect 174954 212058 174986 212614
rect 175542 212058 175574 212614
rect 174954 176614 175574 212058
rect 174954 176058 174986 176614
rect 175542 176058 175574 176614
rect 174954 140614 175574 176058
rect 174954 140058 174986 140614
rect 175542 140058 175574 140614
rect 174954 104614 175574 140058
rect 174954 104058 174986 104614
rect 175542 104058 175574 104614
rect 174954 68614 175574 104058
rect 174954 68058 174986 68614
rect 175542 68058 175574 68614
rect 174954 32614 175574 68058
rect 174954 32058 174986 32614
rect 175542 32058 175574 32614
rect 156954 -6662 156986 -6106
rect 157542 -6662 157574 -6106
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 704838 182414 705830
rect 181794 704282 181826 704838
rect 182382 704282 182414 704838
rect 181794 687454 182414 704282
rect 181794 686898 181826 687454
rect 182382 686898 182414 687454
rect 181794 651454 182414 686898
rect 181794 650898 181826 651454
rect 182382 650898 182414 651454
rect 181794 615454 182414 650898
rect 181794 614898 181826 615454
rect 182382 614898 182414 615454
rect 181794 579454 182414 614898
rect 181794 578898 181826 579454
rect 182382 578898 182414 579454
rect 181794 543454 182414 578898
rect 181794 542898 181826 543454
rect 182382 542898 182414 543454
rect 181794 507454 182414 542898
rect 181794 506898 181826 507454
rect 182382 506898 182414 507454
rect 181794 471454 182414 506898
rect 181794 470898 181826 471454
rect 182382 470898 182414 471454
rect 181794 435454 182414 470898
rect 181794 434898 181826 435454
rect 182382 434898 182414 435454
rect 181794 399454 182414 434898
rect 181794 398898 181826 399454
rect 182382 398898 182414 399454
rect 181794 363454 182414 398898
rect 181794 362898 181826 363454
rect 182382 362898 182414 363454
rect 181794 327454 182414 362898
rect 181794 326898 181826 327454
rect 182382 326898 182414 327454
rect 181794 291454 182414 326898
rect 181794 290898 181826 291454
rect 182382 290898 182414 291454
rect 181794 255454 182414 290898
rect 181794 254898 181826 255454
rect 182382 254898 182414 255454
rect 181794 219454 182414 254898
rect 181794 218898 181826 219454
rect 182382 218898 182414 219454
rect 181794 183454 182414 218898
rect 181794 182898 181826 183454
rect 182382 182898 182414 183454
rect 181794 147454 182414 182898
rect 181794 146898 181826 147454
rect 182382 146898 182414 147454
rect 181794 111454 182414 146898
rect 181794 110898 181826 111454
rect 182382 110898 182414 111454
rect 181794 75454 182414 110898
rect 181794 74898 181826 75454
rect 182382 74898 182414 75454
rect 181794 39454 182414 74898
rect 181794 38898 181826 39454
rect 182382 38898 182414 39454
rect 181794 3454 182414 38898
rect 181794 2898 181826 3454
rect 182382 2898 182414 3454
rect 181794 -346 182414 2898
rect 181794 -902 181826 -346
rect 182382 -902 182414 -346
rect 181794 -1894 182414 -902
rect 185514 691174 186134 706202
rect 185514 690618 185546 691174
rect 186102 690618 186134 691174
rect 185514 655174 186134 690618
rect 185514 654618 185546 655174
rect 186102 654618 186134 655174
rect 185514 619174 186134 654618
rect 185514 618618 185546 619174
rect 186102 618618 186134 619174
rect 185514 583174 186134 618618
rect 185514 582618 185546 583174
rect 186102 582618 186134 583174
rect 185514 547174 186134 582618
rect 185514 546618 185546 547174
rect 186102 546618 186134 547174
rect 185514 511174 186134 546618
rect 185514 510618 185546 511174
rect 186102 510618 186134 511174
rect 185514 475174 186134 510618
rect 185514 474618 185546 475174
rect 186102 474618 186134 475174
rect 185514 439174 186134 474618
rect 185514 438618 185546 439174
rect 186102 438618 186134 439174
rect 185514 403174 186134 438618
rect 185514 402618 185546 403174
rect 186102 402618 186134 403174
rect 185514 367174 186134 402618
rect 185514 366618 185546 367174
rect 186102 366618 186134 367174
rect 185514 331174 186134 366618
rect 185514 330618 185546 331174
rect 186102 330618 186134 331174
rect 185514 295174 186134 330618
rect 185514 294618 185546 295174
rect 186102 294618 186134 295174
rect 185514 259174 186134 294618
rect 185514 258618 185546 259174
rect 186102 258618 186134 259174
rect 185514 223174 186134 258618
rect 185514 222618 185546 223174
rect 186102 222618 186134 223174
rect 185514 187174 186134 222618
rect 185514 186618 185546 187174
rect 186102 186618 186134 187174
rect 185514 151174 186134 186618
rect 185514 150618 185546 151174
rect 186102 150618 186134 151174
rect 185514 115174 186134 150618
rect 185514 114618 185546 115174
rect 186102 114618 186134 115174
rect 185514 79174 186134 114618
rect 185514 78618 185546 79174
rect 186102 78618 186134 79174
rect 185514 43174 186134 78618
rect 185514 42618 185546 43174
rect 186102 42618 186134 43174
rect 185514 7174 186134 42618
rect 185514 6618 185546 7174
rect 186102 6618 186134 7174
rect 185514 -2266 186134 6618
rect 185514 -2822 185546 -2266
rect 186102 -2822 186134 -2266
rect 185514 -3814 186134 -2822
rect 189234 694894 189854 708122
rect 189234 694338 189266 694894
rect 189822 694338 189854 694894
rect 189234 658894 189854 694338
rect 189234 658338 189266 658894
rect 189822 658338 189854 658894
rect 189234 622894 189854 658338
rect 189234 622338 189266 622894
rect 189822 622338 189854 622894
rect 189234 586894 189854 622338
rect 189234 586338 189266 586894
rect 189822 586338 189854 586894
rect 189234 550894 189854 586338
rect 189234 550338 189266 550894
rect 189822 550338 189854 550894
rect 189234 514894 189854 550338
rect 189234 514338 189266 514894
rect 189822 514338 189854 514894
rect 189234 478894 189854 514338
rect 189234 478338 189266 478894
rect 189822 478338 189854 478894
rect 189234 442894 189854 478338
rect 189234 442338 189266 442894
rect 189822 442338 189854 442894
rect 189234 406894 189854 442338
rect 189234 406338 189266 406894
rect 189822 406338 189854 406894
rect 189234 370894 189854 406338
rect 189234 370338 189266 370894
rect 189822 370338 189854 370894
rect 189234 334894 189854 370338
rect 189234 334338 189266 334894
rect 189822 334338 189854 334894
rect 189234 298894 189854 334338
rect 189234 298338 189266 298894
rect 189822 298338 189854 298894
rect 189234 262894 189854 298338
rect 189234 262338 189266 262894
rect 189822 262338 189854 262894
rect 189234 226894 189854 262338
rect 189234 226338 189266 226894
rect 189822 226338 189854 226894
rect 189234 190894 189854 226338
rect 189234 190338 189266 190894
rect 189822 190338 189854 190894
rect 189234 154894 189854 190338
rect 189234 154338 189266 154894
rect 189822 154338 189854 154894
rect 189234 118894 189854 154338
rect 189234 118338 189266 118894
rect 189822 118338 189854 118894
rect 189234 82894 189854 118338
rect 189234 82338 189266 82894
rect 189822 82338 189854 82894
rect 189234 46894 189854 82338
rect 189234 46338 189266 46894
rect 189822 46338 189854 46894
rect 189234 10894 189854 46338
rect 189234 10338 189266 10894
rect 189822 10338 189854 10894
rect 189234 -4186 189854 10338
rect 189234 -4742 189266 -4186
rect 189822 -4742 189854 -4186
rect 189234 -5734 189854 -4742
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711002 210986 711558
rect 211542 711002 211574 711558
rect 207234 709638 207854 709670
rect 207234 709082 207266 709638
rect 207822 709082 207854 709638
rect 203514 707718 204134 707750
rect 203514 707162 203546 707718
rect 204102 707162 204134 707718
rect 192954 698058 192986 698614
rect 193542 698058 193574 698614
rect 192954 662614 193574 698058
rect 192954 662058 192986 662614
rect 193542 662058 193574 662614
rect 192954 626614 193574 662058
rect 192954 626058 192986 626614
rect 193542 626058 193574 626614
rect 192954 590614 193574 626058
rect 192954 590058 192986 590614
rect 193542 590058 193574 590614
rect 192954 554614 193574 590058
rect 192954 554058 192986 554614
rect 193542 554058 193574 554614
rect 192954 518614 193574 554058
rect 192954 518058 192986 518614
rect 193542 518058 193574 518614
rect 192954 482614 193574 518058
rect 192954 482058 192986 482614
rect 193542 482058 193574 482614
rect 192954 446614 193574 482058
rect 192954 446058 192986 446614
rect 193542 446058 193574 446614
rect 192954 410614 193574 446058
rect 192954 410058 192986 410614
rect 193542 410058 193574 410614
rect 192954 374614 193574 410058
rect 192954 374058 192986 374614
rect 193542 374058 193574 374614
rect 192954 338614 193574 374058
rect 192954 338058 192986 338614
rect 193542 338058 193574 338614
rect 192954 302614 193574 338058
rect 192954 302058 192986 302614
rect 193542 302058 193574 302614
rect 192954 266614 193574 302058
rect 192954 266058 192986 266614
rect 193542 266058 193574 266614
rect 192954 230614 193574 266058
rect 192954 230058 192986 230614
rect 193542 230058 193574 230614
rect 192954 194614 193574 230058
rect 192954 194058 192986 194614
rect 193542 194058 193574 194614
rect 192954 158614 193574 194058
rect 192954 158058 192986 158614
rect 193542 158058 193574 158614
rect 192954 122614 193574 158058
rect 192954 122058 192986 122614
rect 193542 122058 193574 122614
rect 192954 86614 193574 122058
rect 192954 86058 192986 86614
rect 193542 86058 193574 86614
rect 192954 50614 193574 86058
rect 192954 50058 192986 50614
rect 193542 50058 193574 50614
rect 192954 14614 193574 50058
rect 192954 14058 192986 14614
rect 193542 14058 193574 14614
rect 174954 -7622 174986 -7066
rect 175542 -7622 175574 -7066
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 705798 200414 705830
rect 199794 705242 199826 705798
rect 200382 705242 200414 705798
rect 199794 669454 200414 705242
rect 199794 668898 199826 669454
rect 200382 668898 200414 669454
rect 199794 633454 200414 668898
rect 199794 632898 199826 633454
rect 200382 632898 200414 633454
rect 199794 597454 200414 632898
rect 199794 596898 199826 597454
rect 200382 596898 200414 597454
rect 199794 561454 200414 596898
rect 199794 560898 199826 561454
rect 200382 560898 200414 561454
rect 199794 525454 200414 560898
rect 199794 524898 199826 525454
rect 200382 524898 200414 525454
rect 199794 489454 200414 524898
rect 199794 488898 199826 489454
rect 200382 488898 200414 489454
rect 199794 453454 200414 488898
rect 199794 452898 199826 453454
rect 200382 452898 200414 453454
rect 199794 417454 200414 452898
rect 199794 416898 199826 417454
rect 200382 416898 200414 417454
rect 199794 381454 200414 416898
rect 199794 380898 199826 381454
rect 200382 380898 200414 381454
rect 199794 345454 200414 380898
rect 199794 344898 199826 345454
rect 200382 344898 200414 345454
rect 199794 309454 200414 344898
rect 199794 308898 199826 309454
rect 200382 308898 200414 309454
rect 199794 273454 200414 308898
rect 199794 272898 199826 273454
rect 200382 272898 200414 273454
rect 199794 237454 200414 272898
rect 199794 236898 199826 237454
rect 200382 236898 200414 237454
rect 199794 201454 200414 236898
rect 199794 200898 199826 201454
rect 200382 200898 200414 201454
rect 199794 165454 200414 200898
rect 199794 164898 199826 165454
rect 200382 164898 200414 165454
rect 199794 129454 200414 164898
rect 199794 128898 199826 129454
rect 200382 128898 200414 129454
rect 199794 93454 200414 128898
rect 199794 92898 199826 93454
rect 200382 92898 200414 93454
rect 199794 57454 200414 92898
rect 199794 56898 199826 57454
rect 200382 56898 200414 57454
rect 199794 21454 200414 56898
rect 199794 20898 199826 21454
rect 200382 20898 200414 21454
rect 199794 -1306 200414 20898
rect 199794 -1862 199826 -1306
rect 200382 -1862 200414 -1306
rect 199794 -1894 200414 -1862
rect 203514 673174 204134 707162
rect 203514 672618 203546 673174
rect 204102 672618 204134 673174
rect 203514 637174 204134 672618
rect 203514 636618 203546 637174
rect 204102 636618 204134 637174
rect 203514 601174 204134 636618
rect 203514 600618 203546 601174
rect 204102 600618 204134 601174
rect 203514 565174 204134 600618
rect 203514 564618 203546 565174
rect 204102 564618 204134 565174
rect 203514 529174 204134 564618
rect 203514 528618 203546 529174
rect 204102 528618 204134 529174
rect 203514 493174 204134 528618
rect 203514 492618 203546 493174
rect 204102 492618 204134 493174
rect 203514 457174 204134 492618
rect 203514 456618 203546 457174
rect 204102 456618 204134 457174
rect 203514 421174 204134 456618
rect 203514 420618 203546 421174
rect 204102 420618 204134 421174
rect 203514 385174 204134 420618
rect 203514 384618 203546 385174
rect 204102 384618 204134 385174
rect 203514 349174 204134 384618
rect 203514 348618 203546 349174
rect 204102 348618 204134 349174
rect 203514 313174 204134 348618
rect 203514 312618 203546 313174
rect 204102 312618 204134 313174
rect 203514 277174 204134 312618
rect 203514 276618 203546 277174
rect 204102 276618 204134 277174
rect 203514 241174 204134 276618
rect 203514 240618 203546 241174
rect 204102 240618 204134 241174
rect 203514 205174 204134 240618
rect 203514 204618 203546 205174
rect 204102 204618 204134 205174
rect 203514 169174 204134 204618
rect 203514 168618 203546 169174
rect 204102 168618 204134 169174
rect 203514 133174 204134 168618
rect 203514 132618 203546 133174
rect 204102 132618 204134 133174
rect 203514 97174 204134 132618
rect 203514 96618 203546 97174
rect 204102 96618 204134 97174
rect 203514 61174 204134 96618
rect 203514 60618 203546 61174
rect 204102 60618 204134 61174
rect 203514 25174 204134 60618
rect 203514 24618 203546 25174
rect 204102 24618 204134 25174
rect 203514 -3226 204134 24618
rect 203514 -3782 203546 -3226
rect 204102 -3782 204134 -3226
rect 203514 -3814 204134 -3782
rect 207234 676894 207854 709082
rect 207234 676338 207266 676894
rect 207822 676338 207854 676894
rect 207234 640894 207854 676338
rect 207234 640338 207266 640894
rect 207822 640338 207854 640894
rect 207234 604894 207854 640338
rect 207234 604338 207266 604894
rect 207822 604338 207854 604894
rect 207234 568894 207854 604338
rect 207234 568338 207266 568894
rect 207822 568338 207854 568894
rect 207234 532894 207854 568338
rect 207234 532338 207266 532894
rect 207822 532338 207854 532894
rect 207234 496894 207854 532338
rect 207234 496338 207266 496894
rect 207822 496338 207854 496894
rect 207234 460894 207854 496338
rect 207234 460338 207266 460894
rect 207822 460338 207854 460894
rect 207234 424894 207854 460338
rect 207234 424338 207266 424894
rect 207822 424338 207854 424894
rect 207234 388894 207854 424338
rect 207234 388338 207266 388894
rect 207822 388338 207854 388894
rect 207234 352894 207854 388338
rect 207234 352338 207266 352894
rect 207822 352338 207854 352894
rect 207234 316894 207854 352338
rect 207234 316338 207266 316894
rect 207822 316338 207854 316894
rect 207234 280894 207854 316338
rect 207234 280338 207266 280894
rect 207822 280338 207854 280894
rect 207234 244894 207854 280338
rect 207234 244338 207266 244894
rect 207822 244338 207854 244894
rect 207234 208894 207854 244338
rect 207234 208338 207266 208894
rect 207822 208338 207854 208894
rect 207234 172894 207854 208338
rect 207234 172338 207266 172894
rect 207822 172338 207854 172894
rect 207234 136894 207854 172338
rect 207234 136338 207266 136894
rect 207822 136338 207854 136894
rect 207234 100894 207854 136338
rect 207234 100338 207266 100894
rect 207822 100338 207854 100894
rect 207234 64894 207854 100338
rect 207234 64338 207266 64894
rect 207822 64338 207854 64894
rect 207234 28894 207854 64338
rect 207234 28338 207266 28894
rect 207822 28338 207854 28894
rect 207234 -5146 207854 28338
rect 207234 -5702 207266 -5146
rect 207822 -5702 207854 -5146
rect 207234 -5734 207854 -5702
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710042 228986 710598
rect 229542 710042 229574 710598
rect 225234 708678 225854 709670
rect 225234 708122 225266 708678
rect 225822 708122 225854 708678
rect 221514 706758 222134 707750
rect 221514 706202 221546 706758
rect 222102 706202 222134 706758
rect 210954 680058 210986 680614
rect 211542 680058 211574 680614
rect 210954 644614 211574 680058
rect 210954 644058 210986 644614
rect 211542 644058 211574 644614
rect 210954 608614 211574 644058
rect 210954 608058 210986 608614
rect 211542 608058 211574 608614
rect 210954 572614 211574 608058
rect 210954 572058 210986 572614
rect 211542 572058 211574 572614
rect 210954 536614 211574 572058
rect 210954 536058 210986 536614
rect 211542 536058 211574 536614
rect 210954 500614 211574 536058
rect 210954 500058 210986 500614
rect 211542 500058 211574 500614
rect 210954 464614 211574 500058
rect 210954 464058 210986 464614
rect 211542 464058 211574 464614
rect 210954 428614 211574 464058
rect 210954 428058 210986 428614
rect 211542 428058 211574 428614
rect 210954 392614 211574 428058
rect 210954 392058 210986 392614
rect 211542 392058 211574 392614
rect 210954 356614 211574 392058
rect 210954 356058 210986 356614
rect 211542 356058 211574 356614
rect 210954 320614 211574 356058
rect 210954 320058 210986 320614
rect 211542 320058 211574 320614
rect 210954 284614 211574 320058
rect 210954 284058 210986 284614
rect 211542 284058 211574 284614
rect 210954 248614 211574 284058
rect 210954 248058 210986 248614
rect 211542 248058 211574 248614
rect 210954 212614 211574 248058
rect 210954 212058 210986 212614
rect 211542 212058 211574 212614
rect 210954 176614 211574 212058
rect 210954 176058 210986 176614
rect 211542 176058 211574 176614
rect 210954 140614 211574 176058
rect 210954 140058 210986 140614
rect 211542 140058 211574 140614
rect 210954 104614 211574 140058
rect 210954 104058 210986 104614
rect 211542 104058 211574 104614
rect 210954 68614 211574 104058
rect 210954 68058 210986 68614
rect 211542 68058 211574 68614
rect 210954 32614 211574 68058
rect 210954 32058 210986 32614
rect 211542 32058 211574 32614
rect 192954 -6662 192986 -6106
rect 193542 -6662 193574 -6106
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 704838 218414 705830
rect 217794 704282 217826 704838
rect 218382 704282 218414 704838
rect 217794 687454 218414 704282
rect 217794 686898 217826 687454
rect 218382 686898 218414 687454
rect 217794 651454 218414 686898
rect 217794 650898 217826 651454
rect 218382 650898 218414 651454
rect 217794 615454 218414 650898
rect 217794 614898 217826 615454
rect 218382 614898 218414 615454
rect 217794 579454 218414 614898
rect 217794 578898 217826 579454
rect 218382 578898 218414 579454
rect 217794 543454 218414 578898
rect 217794 542898 217826 543454
rect 218382 542898 218414 543454
rect 217794 507454 218414 542898
rect 217794 506898 217826 507454
rect 218382 506898 218414 507454
rect 217794 471454 218414 506898
rect 217794 470898 217826 471454
rect 218382 470898 218414 471454
rect 217794 435454 218414 470898
rect 217794 434898 217826 435454
rect 218382 434898 218414 435454
rect 217794 399454 218414 434898
rect 217794 398898 217826 399454
rect 218382 398898 218414 399454
rect 217794 363454 218414 398898
rect 217794 362898 217826 363454
rect 218382 362898 218414 363454
rect 217794 327454 218414 362898
rect 217794 326898 217826 327454
rect 218382 326898 218414 327454
rect 217794 291454 218414 326898
rect 217794 290898 217826 291454
rect 218382 290898 218414 291454
rect 217794 255454 218414 290898
rect 217794 254898 217826 255454
rect 218382 254898 218414 255454
rect 217794 219454 218414 254898
rect 217794 218898 217826 219454
rect 218382 218898 218414 219454
rect 217794 183454 218414 218898
rect 217794 182898 217826 183454
rect 218382 182898 218414 183454
rect 217794 147454 218414 182898
rect 217794 146898 217826 147454
rect 218382 146898 218414 147454
rect 217794 111454 218414 146898
rect 217794 110898 217826 111454
rect 218382 110898 218414 111454
rect 217794 75454 218414 110898
rect 217794 74898 217826 75454
rect 218382 74898 218414 75454
rect 217794 39454 218414 74898
rect 217794 38898 217826 39454
rect 218382 38898 218414 39454
rect 217794 3454 218414 38898
rect 217794 2898 217826 3454
rect 218382 2898 218414 3454
rect 217794 -346 218414 2898
rect 217794 -902 217826 -346
rect 218382 -902 218414 -346
rect 217794 -1894 218414 -902
rect 221514 691174 222134 706202
rect 221514 690618 221546 691174
rect 222102 690618 222134 691174
rect 221514 655174 222134 690618
rect 221514 654618 221546 655174
rect 222102 654618 222134 655174
rect 221514 619174 222134 654618
rect 221514 618618 221546 619174
rect 222102 618618 222134 619174
rect 221514 583174 222134 618618
rect 221514 582618 221546 583174
rect 222102 582618 222134 583174
rect 221514 547174 222134 582618
rect 221514 546618 221546 547174
rect 222102 546618 222134 547174
rect 221514 511174 222134 546618
rect 221514 510618 221546 511174
rect 222102 510618 222134 511174
rect 221514 475174 222134 510618
rect 221514 474618 221546 475174
rect 222102 474618 222134 475174
rect 221514 439174 222134 474618
rect 221514 438618 221546 439174
rect 222102 438618 222134 439174
rect 221514 403174 222134 438618
rect 221514 402618 221546 403174
rect 222102 402618 222134 403174
rect 221514 367174 222134 402618
rect 221514 366618 221546 367174
rect 222102 366618 222134 367174
rect 221514 331174 222134 366618
rect 221514 330618 221546 331174
rect 222102 330618 222134 331174
rect 221514 295174 222134 330618
rect 221514 294618 221546 295174
rect 222102 294618 222134 295174
rect 221514 259174 222134 294618
rect 221514 258618 221546 259174
rect 222102 258618 222134 259174
rect 221514 223174 222134 258618
rect 221514 222618 221546 223174
rect 222102 222618 222134 223174
rect 221514 187174 222134 222618
rect 221514 186618 221546 187174
rect 222102 186618 222134 187174
rect 221514 151174 222134 186618
rect 221514 150618 221546 151174
rect 222102 150618 222134 151174
rect 221514 115174 222134 150618
rect 221514 114618 221546 115174
rect 222102 114618 222134 115174
rect 221514 79174 222134 114618
rect 221514 78618 221546 79174
rect 222102 78618 222134 79174
rect 221514 43174 222134 78618
rect 221514 42618 221546 43174
rect 222102 42618 222134 43174
rect 221514 7174 222134 42618
rect 221514 6618 221546 7174
rect 222102 6618 222134 7174
rect 221514 -2266 222134 6618
rect 221514 -2822 221546 -2266
rect 222102 -2822 222134 -2266
rect 221514 -3814 222134 -2822
rect 225234 694894 225854 708122
rect 225234 694338 225266 694894
rect 225822 694338 225854 694894
rect 225234 658894 225854 694338
rect 225234 658338 225266 658894
rect 225822 658338 225854 658894
rect 225234 622894 225854 658338
rect 225234 622338 225266 622894
rect 225822 622338 225854 622894
rect 225234 586894 225854 622338
rect 225234 586338 225266 586894
rect 225822 586338 225854 586894
rect 225234 550894 225854 586338
rect 225234 550338 225266 550894
rect 225822 550338 225854 550894
rect 225234 514894 225854 550338
rect 225234 514338 225266 514894
rect 225822 514338 225854 514894
rect 225234 478894 225854 514338
rect 225234 478338 225266 478894
rect 225822 478338 225854 478894
rect 225234 442894 225854 478338
rect 225234 442338 225266 442894
rect 225822 442338 225854 442894
rect 225234 406894 225854 442338
rect 225234 406338 225266 406894
rect 225822 406338 225854 406894
rect 225234 370894 225854 406338
rect 225234 370338 225266 370894
rect 225822 370338 225854 370894
rect 225234 334894 225854 370338
rect 225234 334338 225266 334894
rect 225822 334338 225854 334894
rect 225234 298894 225854 334338
rect 225234 298338 225266 298894
rect 225822 298338 225854 298894
rect 225234 262894 225854 298338
rect 225234 262338 225266 262894
rect 225822 262338 225854 262894
rect 225234 226894 225854 262338
rect 225234 226338 225266 226894
rect 225822 226338 225854 226894
rect 225234 190894 225854 226338
rect 225234 190338 225266 190894
rect 225822 190338 225854 190894
rect 225234 154894 225854 190338
rect 225234 154338 225266 154894
rect 225822 154338 225854 154894
rect 225234 118894 225854 154338
rect 225234 118338 225266 118894
rect 225822 118338 225854 118894
rect 225234 82894 225854 118338
rect 225234 82338 225266 82894
rect 225822 82338 225854 82894
rect 225234 46894 225854 82338
rect 225234 46338 225266 46894
rect 225822 46338 225854 46894
rect 225234 10894 225854 46338
rect 225234 10338 225266 10894
rect 225822 10338 225854 10894
rect 225234 -4186 225854 10338
rect 225234 -4742 225266 -4186
rect 225822 -4742 225854 -4186
rect 225234 -5734 225854 -4742
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711002 246986 711558
rect 247542 711002 247574 711558
rect 243234 709638 243854 709670
rect 243234 709082 243266 709638
rect 243822 709082 243854 709638
rect 239514 707718 240134 707750
rect 239514 707162 239546 707718
rect 240102 707162 240134 707718
rect 228954 698058 228986 698614
rect 229542 698058 229574 698614
rect 228954 662614 229574 698058
rect 228954 662058 228986 662614
rect 229542 662058 229574 662614
rect 228954 626614 229574 662058
rect 228954 626058 228986 626614
rect 229542 626058 229574 626614
rect 228954 590614 229574 626058
rect 228954 590058 228986 590614
rect 229542 590058 229574 590614
rect 228954 554614 229574 590058
rect 228954 554058 228986 554614
rect 229542 554058 229574 554614
rect 228954 518614 229574 554058
rect 228954 518058 228986 518614
rect 229542 518058 229574 518614
rect 228954 482614 229574 518058
rect 228954 482058 228986 482614
rect 229542 482058 229574 482614
rect 228954 446614 229574 482058
rect 235794 705798 236414 705830
rect 235794 705242 235826 705798
rect 236382 705242 236414 705798
rect 235794 669454 236414 705242
rect 235794 668898 235826 669454
rect 236382 668898 236414 669454
rect 235794 633454 236414 668898
rect 235794 632898 235826 633454
rect 236382 632898 236414 633454
rect 235794 597454 236414 632898
rect 235794 596898 235826 597454
rect 236382 596898 236414 597454
rect 235794 561454 236414 596898
rect 235794 560898 235826 561454
rect 236382 560898 236414 561454
rect 235794 525454 236414 560898
rect 235794 524898 235826 525454
rect 236382 524898 236414 525454
rect 235794 489454 236414 524898
rect 235794 488898 235826 489454
rect 236382 488898 236414 489454
rect 235794 458000 236414 488898
rect 239514 673174 240134 707162
rect 239514 672618 239546 673174
rect 240102 672618 240134 673174
rect 239514 637174 240134 672618
rect 239514 636618 239546 637174
rect 240102 636618 240134 637174
rect 239514 601174 240134 636618
rect 239514 600618 239546 601174
rect 240102 600618 240134 601174
rect 239514 565174 240134 600618
rect 239514 564618 239546 565174
rect 240102 564618 240134 565174
rect 239514 529174 240134 564618
rect 239514 528618 239546 529174
rect 240102 528618 240134 529174
rect 239514 493174 240134 528618
rect 239514 492618 239546 493174
rect 240102 492618 240134 493174
rect 239514 460000 240134 492618
rect 243234 676894 243854 709082
rect 243234 676338 243266 676894
rect 243822 676338 243854 676894
rect 243234 640894 243854 676338
rect 243234 640338 243266 640894
rect 243822 640338 243854 640894
rect 243234 604894 243854 640338
rect 243234 604338 243266 604894
rect 243822 604338 243854 604894
rect 243234 568894 243854 604338
rect 243234 568338 243266 568894
rect 243822 568338 243854 568894
rect 243234 532894 243854 568338
rect 243234 532338 243266 532894
rect 243822 532338 243854 532894
rect 243234 496894 243854 532338
rect 243234 496338 243266 496894
rect 243822 496338 243854 496894
rect 243234 460894 243854 496338
rect 243234 460338 243266 460894
rect 243822 460338 243854 460894
rect 243234 460000 243854 460338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710042 264986 710598
rect 265542 710042 265574 710598
rect 261234 708678 261854 709670
rect 261234 708122 261266 708678
rect 261822 708122 261854 708678
rect 257514 706758 258134 707750
rect 257514 706202 257546 706758
rect 258102 706202 258134 706758
rect 246954 680058 246986 680614
rect 247542 680058 247574 680614
rect 246954 644614 247574 680058
rect 246954 644058 246986 644614
rect 247542 644058 247574 644614
rect 246954 608614 247574 644058
rect 246954 608058 246986 608614
rect 247542 608058 247574 608614
rect 246954 572614 247574 608058
rect 246954 572058 246986 572614
rect 247542 572058 247574 572614
rect 246954 536614 247574 572058
rect 246954 536058 246986 536614
rect 247542 536058 247574 536614
rect 246954 500614 247574 536058
rect 246954 500058 246986 500614
rect 247542 500058 247574 500614
rect 246954 464614 247574 500058
rect 246954 464058 246986 464614
rect 247542 464058 247574 464614
rect 246954 460000 247574 464058
rect 253794 704838 254414 705830
rect 253794 704282 253826 704838
rect 254382 704282 254414 704838
rect 253794 687454 254414 704282
rect 253794 686898 253826 687454
rect 254382 686898 254414 687454
rect 253794 651454 254414 686898
rect 253794 650898 253826 651454
rect 254382 650898 254414 651454
rect 253794 615454 254414 650898
rect 253794 614898 253826 615454
rect 254382 614898 254414 615454
rect 253794 579454 254414 614898
rect 253794 578898 253826 579454
rect 254382 578898 254414 579454
rect 253794 543454 254414 578898
rect 253794 542898 253826 543454
rect 254382 542898 254414 543454
rect 253794 507454 254414 542898
rect 253794 506898 253826 507454
rect 254382 506898 254414 507454
rect 253794 471454 254414 506898
rect 253794 470898 253826 471454
rect 254382 470898 254414 471454
rect 253794 458000 254414 470898
rect 257514 691174 258134 706202
rect 257514 690618 257546 691174
rect 258102 690618 258134 691174
rect 257514 655174 258134 690618
rect 257514 654618 257546 655174
rect 258102 654618 258134 655174
rect 257514 619174 258134 654618
rect 257514 618618 257546 619174
rect 258102 618618 258134 619174
rect 257514 583174 258134 618618
rect 257514 582618 257546 583174
rect 258102 582618 258134 583174
rect 257514 547174 258134 582618
rect 257514 546618 257546 547174
rect 258102 546618 258134 547174
rect 257514 511174 258134 546618
rect 257514 510618 257546 511174
rect 258102 510618 258134 511174
rect 257514 475174 258134 510618
rect 257514 474618 257546 475174
rect 258102 474618 258134 475174
rect 257514 460000 258134 474618
rect 261234 694894 261854 708122
rect 261234 694338 261266 694894
rect 261822 694338 261854 694894
rect 261234 658894 261854 694338
rect 261234 658338 261266 658894
rect 261822 658338 261854 658894
rect 261234 622894 261854 658338
rect 261234 622338 261266 622894
rect 261822 622338 261854 622894
rect 261234 586894 261854 622338
rect 261234 586338 261266 586894
rect 261822 586338 261854 586894
rect 261234 550894 261854 586338
rect 261234 550338 261266 550894
rect 261822 550338 261854 550894
rect 261234 514894 261854 550338
rect 261234 514338 261266 514894
rect 261822 514338 261854 514894
rect 261234 478894 261854 514338
rect 261234 478338 261266 478894
rect 261822 478338 261854 478894
rect 261234 460000 261854 478338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711002 282986 711558
rect 283542 711002 283574 711558
rect 279234 709638 279854 709670
rect 279234 709082 279266 709638
rect 279822 709082 279854 709638
rect 275514 707718 276134 707750
rect 275514 707162 275546 707718
rect 276102 707162 276134 707718
rect 264954 698058 264986 698614
rect 265542 698058 265574 698614
rect 264954 662614 265574 698058
rect 264954 662058 264986 662614
rect 265542 662058 265574 662614
rect 264954 626614 265574 662058
rect 264954 626058 264986 626614
rect 265542 626058 265574 626614
rect 264954 590614 265574 626058
rect 264954 590058 264986 590614
rect 265542 590058 265574 590614
rect 264954 554614 265574 590058
rect 264954 554058 264986 554614
rect 265542 554058 265574 554614
rect 264954 518614 265574 554058
rect 264954 518058 264986 518614
rect 265542 518058 265574 518614
rect 264954 482614 265574 518058
rect 264954 482058 264986 482614
rect 265542 482058 265574 482614
rect 264954 460000 265574 482058
rect 271794 705798 272414 705830
rect 271794 705242 271826 705798
rect 272382 705242 272414 705798
rect 271794 669454 272414 705242
rect 271794 668898 271826 669454
rect 272382 668898 272414 669454
rect 271794 633454 272414 668898
rect 271794 632898 271826 633454
rect 272382 632898 272414 633454
rect 271794 597454 272414 632898
rect 271794 596898 271826 597454
rect 272382 596898 272414 597454
rect 271794 561454 272414 596898
rect 271794 560898 271826 561454
rect 272382 560898 272414 561454
rect 271794 525454 272414 560898
rect 271794 524898 271826 525454
rect 272382 524898 272414 525454
rect 271794 489454 272414 524898
rect 271794 488898 271826 489454
rect 272382 488898 272414 489454
rect 271794 458000 272414 488898
rect 275514 673174 276134 707162
rect 275514 672618 275546 673174
rect 276102 672618 276134 673174
rect 275514 637174 276134 672618
rect 275514 636618 275546 637174
rect 276102 636618 276134 637174
rect 275514 601174 276134 636618
rect 275514 600618 275546 601174
rect 276102 600618 276134 601174
rect 275514 565174 276134 600618
rect 275514 564618 275546 565174
rect 276102 564618 276134 565174
rect 275514 529174 276134 564618
rect 275514 528618 275546 529174
rect 276102 528618 276134 529174
rect 275514 493174 276134 528618
rect 275514 492618 275546 493174
rect 276102 492618 276134 493174
rect 275514 460000 276134 492618
rect 279234 676894 279854 709082
rect 279234 676338 279266 676894
rect 279822 676338 279854 676894
rect 279234 640894 279854 676338
rect 279234 640338 279266 640894
rect 279822 640338 279854 640894
rect 279234 604894 279854 640338
rect 279234 604338 279266 604894
rect 279822 604338 279854 604894
rect 279234 568894 279854 604338
rect 279234 568338 279266 568894
rect 279822 568338 279854 568894
rect 279234 532894 279854 568338
rect 279234 532338 279266 532894
rect 279822 532338 279854 532894
rect 279234 496894 279854 532338
rect 279234 496338 279266 496894
rect 279822 496338 279854 496894
rect 279234 460894 279854 496338
rect 279234 460338 279266 460894
rect 279822 460338 279854 460894
rect 279234 460000 279854 460338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710042 300986 710598
rect 301542 710042 301574 710598
rect 297234 708678 297854 709670
rect 297234 708122 297266 708678
rect 297822 708122 297854 708678
rect 293514 706758 294134 707750
rect 293514 706202 293546 706758
rect 294102 706202 294134 706758
rect 282954 680058 282986 680614
rect 283542 680058 283574 680614
rect 282954 644614 283574 680058
rect 282954 644058 282986 644614
rect 283542 644058 283574 644614
rect 282954 608614 283574 644058
rect 282954 608058 282986 608614
rect 283542 608058 283574 608614
rect 282954 572614 283574 608058
rect 282954 572058 282986 572614
rect 283542 572058 283574 572614
rect 282954 536614 283574 572058
rect 282954 536058 282986 536614
rect 283542 536058 283574 536614
rect 282954 500614 283574 536058
rect 282954 500058 282986 500614
rect 283542 500058 283574 500614
rect 282954 464614 283574 500058
rect 282954 464058 282986 464614
rect 283542 464058 283574 464614
rect 282954 460000 283574 464058
rect 289794 704838 290414 705830
rect 289794 704282 289826 704838
rect 290382 704282 290414 704838
rect 289794 687454 290414 704282
rect 289794 686898 289826 687454
rect 290382 686898 290414 687454
rect 289794 651454 290414 686898
rect 289794 650898 289826 651454
rect 290382 650898 290414 651454
rect 289794 615454 290414 650898
rect 289794 614898 289826 615454
rect 290382 614898 290414 615454
rect 289794 579454 290414 614898
rect 289794 578898 289826 579454
rect 290382 578898 290414 579454
rect 289794 543454 290414 578898
rect 289794 542898 289826 543454
rect 290382 542898 290414 543454
rect 289794 507454 290414 542898
rect 289794 506898 289826 507454
rect 290382 506898 290414 507454
rect 289794 471454 290414 506898
rect 289794 470898 289826 471454
rect 290382 470898 290414 471454
rect 289794 458000 290414 470898
rect 293514 691174 294134 706202
rect 293514 690618 293546 691174
rect 294102 690618 294134 691174
rect 293514 655174 294134 690618
rect 293514 654618 293546 655174
rect 294102 654618 294134 655174
rect 293514 619174 294134 654618
rect 293514 618618 293546 619174
rect 294102 618618 294134 619174
rect 293514 583174 294134 618618
rect 293514 582618 293546 583174
rect 294102 582618 294134 583174
rect 293514 547174 294134 582618
rect 293514 546618 293546 547174
rect 294102 546618 294134 547174
rect 293514 511174 294134 546618
rect 293514 510618 293546 511174
rect 294102 510618 294134 511174
rect 293514 475174 294134 510618
rect 293514 474618 293546 475174
rect 294102 474618 294134 475174
rect 293514 460000 294134 474618
rect 297234 694894 297854 708122
rect 297234 694338 297266 694894
rect 297822 694338 297854 694894
rect 297234 658894 297854 694338
rect 297234 658338 297266 658894
rect 297822 658338 297854 658894
rect 297234 622894 297854 658338
rect 297234 622338 297266 622894
rect 297822 622338 297854 622894
rect 297234 586894 297854 622338
rect 297234 586338 297266 586894
rect 297822 586338 297854 586894
rect 297234 550894 297854 586338
rect 297234 550338 297266 550894
rect 297822 550338 297854 550894
rect 297234 514894 297854 550338
rect 297234 514338 297266 514894
rect 297822 514338 297854 514894
rect 297234 478894 297854 514338
rect 297234 478338 297266 478894
rect 297822 478338 297854 478894
rect 297234 460000 297854 478338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711002 318986 711558
rect 319542 711002 319574 711558
rect 315234 709638 315854 709670
rect 315234 709082 315266 709638
rect 315822 709082 315854 709638
rect 311514 707718 312134 707750
rect 311514 707162 311546 707718
rect 312102 707162 312134 707718
rect 300954 698058 300986 698614
rect 301542 698058 301574 698614
rect 300954 662614 301574 698058
rect 300954 662058 300986 662614
rect 301542 662058 301574 662614
rect 300954 626614 301574 662058
rect 300954 626058 300986 626614
rect 301542 626058 301574 626614
rect 300954 590614 301574 626058
rect 300954 590058 300986 590614
rect 301542 590058 301574 590614
rect 300954 554614 301574 590058
rect 300954 554058 300986 554614
rect 301542 554058 301574 554614
rect 300954 518614 301574 554058
rect 300954 518058 300986 518614
rect 301542 518058 301574 518614
rect 300954 482614 301574 518058
rect 300954 482058 300986 482614
rect 301542 482058 301574 482614
rect 300954 460000 301574 482058
rect 307794 705798 308414 705830
rect 307794 705242 307826 705798
rect 308382 705242 308414 705798
rect 307794 669454 308414 705242
rect 307794 668898 307826 669454
rect 308382 668898 308414 669454
rect 307794 633454 308414 668898
rect 307794 632898 307826 633454
rect 308382 632898 308414 633454
rect 307794 597454 308414 632898
rect 307794 596898 307826 597454
rect 308382 596898 308414 597454
rect 307794 561454 308414 596898
rect 307794 560898 307826 561454
rect 308382 560898 308414 561454
rect 307794 525454 308414 560898
rect 307794 524898 307826 525454
rect 308382 524898 308414 525454
rect 307794 489454 308414 524898
rect 307794 488898 307826 489454
rect 308382 488898 308414 489454
rect 307794 458000 308414 488898
rect 311514 673174 312134 707162
rect 311514 672618 311546 673174
rect 312102 672618 312134 673174
rect 311514 637174 312134 672618
rect 311514 636618 311546 637174
rect 312102 636618 312134 637174
rect 311514 601174 312134 636618
rect 311514 600618 311546 601174
rect 312102 600618 312134 601174
rect 311514 565174 312134 600618
rect 311514 564618 311546 565174
rect 312102 564618 312134 565174
rect 311514 529174 312134 564618
rect 311514 528618 311546 529174
rect 312102 528618 312134 529174
rect 311514 493174 312134 528618
rect 311514 492618 311546 493174
rect 312102 492618 312134 493174
rect 311514 460000 312134 492618
rect 315234 676894 315854 709082
rect 315234 676338 315266 676894
rect 315822 676338 315854 676894
rect 315234 640894 315854 676338
rect 315234 640338 315266 640894
rect 315822 640338 315854 640894
rect 315234 604894 315854 640338
rect 315234 604338 315266 604894
rect 315822 604338 315854 604894
rect 315234 568894 315854 604338
rect 315234 568338 315266 568894
rect 315822 568338 315854 568894
rect 315234 532894 315854 568338
rect 315234 532338 315266 532894
rect 315822 532338 315854 532894
rect 315234 496894 315854 532338
rect 315234 496338 315266 496894
rect 315822 496338 315854 496894
rect 315234 460894 315854 496338
rect 315234 460338 315266 460894
rect 315822 460338 315854 460894
rect 315234 460000 315854 460338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710042 336986 710598
rect 337542 710042 337574 710598
rect 333234 708678 333854 709670
rect 333234 708122 333266 708678
rect 333822 708122 333854 708678
rect 329514 706758 330134 707750
rect 329514 706202 329546 706758
rect 330102 706202 330134 706758
rect 318954 680058 318986 680614
rect 319542 680058 319574 680614
rect 318954 644614 319574 680058
rect 318954 644058 318986 644614
rect 319542 644058 319574 644614
rect 318954 608614 319574 644058
rect 318954 608058 318986 608614
rect 319542 608058 319574 608614
rect 318954 572614 319574 608058
rect 318954 572058 318986 572614
rect 319542 572058 319574 572614
rect 318954 536614 319574 572058
rect 318954 536058 318986 536614
rect 319542 536058 319574 536614
rect 318954 500614 319574 536058
rect 318954 500058 318986 500614
rect 319542 500058 319574 500614
rect 318954 464614 319574 500058
rect 318954 464058 318986 464614
rect 319542 464058 319574 464614
rect 318954 460000 319574 464058
rect 325794 704838 326414 705830
rect 325794 704282 325826 704838
rect 326382 704282 326414 704838
rect 325794 687454 326414 704282
rect 325794 686898 325826 687454
rect 326382 686898 326414 687454
rect 325794 651454 326414 686898
rect 325794 650898 325826 651454
rect 326382 650898 326414 651454
rect 325794 615454 326414 650898
rect 325794 614898 325826 615454
rect 326382 614898 326414 615454
rect 325794 579454 326414 614898
rect 325794 578898 325826 579454
rect 326382 578898 326414 579454
rect 325794 543454 326414 578898
rect 325794 542898 325826 543454
rect 326382 542898 326414 543454
rect 325794 507454 326414 542898
rect 325794 506898 325826 507454
rect 326382 506898 326414 507454
rect 325794 471454 326414 506898
rect 325794 470898 325826 471454
rect 326382 470898 326414 471454
rect 325794 458000 326414 470898
rect 329514 691174 330134 706202
rect 329514 690618 329546 691174
rect 330102 690618 330134 691174
rect 329514 655174 330134 690618
rect 329514 654618 329546 655174
rect 330102 654618 330134 655174
rect 329514 619174 330134 654618
rect 329514 618618 329546 619174
rect 330102 618618 330134 619174
rect 329514 583174 330134 618618
rect 329514 582618 329546 583174
rect 330102 582618 330134 583174
rect 329514 547174 330134 582618
rect 329514 546618 329546 547174
rect 330102 546618 330134 547174
rect 329514 511174 330134 546618
rect 329514 510618 329546 511174
rect 330102 510618 330134 511174
rect 329514 475174 330134 510618
rect 329514 474618 329546 475174
rect 330102 474618 330134 475174
rect 329514 460000 330134 474618
rect 333234 694894 333854 708122
rect 333234 694338 333266 694894
rect 333822 694338 333854 694894
rect 333234 658894 333854 694338
rect 333234 658338 333266 658894
rect 333822 658338 333854 658894
rect 333234 622894 333854 658338
rect 333234 622338 333266 622894
rect 333822 622338 333854 622894
rect 333234 586894 333854 622338
rect 333234 586338 333266 586894
rect 333822 586338 333854 586894
rect 333234 550894 333854 586338
rect 333234 550338 333266 550894
rect 333822 550338 333854 550894
rect 333234 514894 333854 550338
rect 333234 514338 333266 514894
rect 333822 514338 333854 514894
rect 333234 478894 333854 514338
rect 333234 478338 333266 478894
rect 333822 478338 333854 478894
rect 333234 460000 333854 478338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711002 354986 711558
rect 355542 711002 355574 711558
rect 351234 709638 351854 709670
rect 351234 709082 351266 709638
rect 351822 709082 351854 709638
rect 347514 707718 348134 707750
rect 347514 707162 347546 707718
rect 348102 707162 348134 707718
rect 336954 698058 336986 698614
rect 337542 698058 337574 698614
rect 336954 662614 337574 698058
rect 336954 662058 336986 662614
rect 337542 662058 337574 662614
rect 336954 626614 337574 662058
rect 336954 626058 336986 626614
rect 337542 626058 337574 626614
rect 336954 590614 337574 626058
rect 336954 590058 336986 590614
rect 337542 590058 337574 590614
rect 336954 554614 337574 590058
rect 336954 554058 336986 554614
rect 337542 554058 337574 554614
rect 336954 518614 337574 554058
rect 336954 518058 336986 518614
rect 337542 518058 337574 518614
rect 336954 482614 337574 518058
rect 336954 482058 336986 482614
rect 337542 482058 337574 482614
rect 336954 460000 337574 482058
rect 343794 705798 344414 705830
rect 343794 705242 343826 705798
rect 344382 705242 344414 705798
rect 343794 669454 344414 705242
rect 343794 668898 343826 669454
rect 344382 668898 344414 669454
rect 343794 633454 344414 668898
rect 343794 632898 343826 633454
rect 344382 632898 344414 633454
rect 343794 597454 344414 632898
rect 343794 596898 343826 597454
rect 344382 596898 344414 597454
rect 343794 561454 344414 596898
rect 343794 560898 343826 561454
rect 344382 560898 344414 561454
rect 343794 525454 344414 560898
rect 343794 524898 343826 525454
rect 344382 524898 344414 525454
rect 343794 489454 344414 524898
rect 343794 488898 343826 489454
rect 344382 488898 344414 489454
rect 343794 458000 344414 488898
rect 347514 673174 348134 707162
rect 347514 672618 347546 673174
rect 348102 672618 348134 673174
rect 347514 637174 348134 672618
rect 347514 636618 347546 637174
rect 348102 636618 348134 637174
rect 347514 601174 348134 636618
rect 347514 600618 347546 601174
rect 348102 600618 348134 601174
rect 347514 565174 348134 600618
rect 347514 564618 347546 565174
rect 348102 564618 348134 565174
rect 347514 529174 348134 564618
rect 347514 528618 347546 529174
rect 348102 528618 348134 529174
rect 347514 493174 348134 528618
rect 347514 492618 347546 493174
rect 348102 492618 348134 493174
rect 347514 460000 348134 492618
rect 351234 676894 351854 709082
rect 351234 676338 351266 676894
rect 351822 676338 351854 676894
rect 351234 640894 351854 676338
rect 351234 640338 351266 640894
rect 351822 640338 351854 640894
rect 351234 604894 351854 640338
rect 351234 604338 351266 604894
rect 351822 604338 351854 604894
rect 351234 568894 351854 604338
rect 351234 568338 351266 568894
rect 351822 568338 351854 568894
rect 351234 532894 351854 568338
rect 351234 532338 351266 532894
rect 351822 532338 351854 532894
rect 351234 496894 351854 532338
rect 351234 496338 351266 496894
rect 351822 496338 351854 496894
rect 351234 460894 351854 496338
rect 351234 460338 351266 460894
rect 351822 460338 351854 460894
rect 351234 460000 351854 460338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710042 372986 710598
rect 373542 710042 373574 710598
rect 369234 708678 369854 709670
rect 369234 708122 369266 708678
rect 369822 708122 369854 708678
rect 365514 706758 366134 707750
rect 365514 706202 365546 706758
rect 366102 706202 366134 706758
rect 354954 680058 354986 680614
rect 355542 680058 355574 680614
rect 354954 644614 355574 680058
rect 354954 644058 354986 644614
rect 355542 644058 355574 644614
rect 354954 608614 355574 644058
rect 354954 608058 354986 608614
rect 355542 608058 355574 608614
rect 354954 572614 355574 608058
rect 354954 572058 354986 572614
rect 355542 572058 355574 572614
rect 354954 536614 355574 572058
rect 354954 536058 354986 536614
rect 355542 536058 355574 536614
rect 354954 500614 355574 536058
rect 354954 500058 354986 500614
rect 355542 500058 355574 500614
rect 354954 464614 355574 500058
rect 354954 464058 354986 464614
rect 355542 464058 355574 464614
rect 354954 460000 355574 464058
rect 361794 704838 362414 705830
rect 361794 704282 361826 704838
rect 362382 704282 362414 704838
rect 361794 687454 362414 704282
rect 361794 686898 361826 687454
rect 362382 686898 362414 687454
rect 361794 651454 362414 686898
rect 361794 650898 361826 651454
rect 362382 650898 362414 651454
rect 361794 615454 362414 650898
rect 361794 614898 361826 615454
rect 362382 614898 362414 615454
rect 361794 579454 362414 614898
rect 361794 578898 361826 579454
rect 362382 578898 362414 579454
rect 361794 543454 362414 578898
rect 361794 542898 361826 543454
rect 362382 542898 362414 543454
rect 361794 507454 362414 542898
rect 361794 506898 361826 507454
rect 362382 506898 362414 507454
rect 361794 471454 362414 506898
rect 361794 470898 361826 471454
rect 362382 470898 362414 471454
rect 361794 458000 362414 470898
rect 365514 691174 366134 706202
rect 365514 690618 365546 691174
rect 366102 690618 366134 691174
rect 365514 655174 366134 690618
rect 365514 654618 365546 655174
rect 366102 654618 366134 655174
rect 365514 619174 366134 654618
rect 365514 618618 365546 619174
rect 366102 618618 366134 619174
rect 365514 583174 366134 618618
rect 365514 582618 365546 583174
rect 366102 582618 366134 583174
rect 365514 547174 366134 582618
rect 365514 546618 365546 547174
rect 366102 546618 366134 547174
rect 365514 511174 366134 546618
rect 365514 510618 365546 511174
rect 366102 510618 366134 511174
rect 365514 475174 366134 510618
rect 365514 474618 365546 475174
rect 366102 474618 366134 475174
rect 365514 460000 366134 474618
rect 369234 694894 369854 708122
rect 369234 694338 369266 694894
rect 369822 694338 369854 694894
rect 369234 658894 369854 694338
rect 369234 658338 369266 658894
rect 369822 658338 369854 658894
rect 369234 622894 369854 658338
rect 369234 622338 369266 622894
rect 369822 622338 369854 622894
rect 369234 586894 369854 622338
rect 369234 586338 369266 586894
rect 369822 586338 369854 586894
rect 369234 550894 369854 586338
rect 369234 550338 369266 550894
rect 369822 550338 369854 550894
rect 369234 514894 369854 550338
rect 369234 514338 369266 514894
rect 369822 514338 369854 514894
rect 369234 478894 369854 514338
rect 369234 478338 369266 478894
rect 369822 478338 369854 478894
rect 369234 460000 369854 478338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711002 390986 711558
rect 391542 711002 391574 711558
rect 387234 709638 387854 709670
rect 387234 709082 387266 709638
rect 387822 709082 387854 709638
rect 383514 707718 384134 707750
rect 383514 707162 383546 707718
rect 384102 707162 384134 707718
rect 372954 698058 372986 698614
rect 373542 698058 373574 698614
rect 372954 662614 373574 698058
rect 372954 662058 372986 662614
rect 373542 662058 373574 662614
rect 372954 626614 373574 662058
rect 372954 626058 372986 626614
rect 373542 626058 373574 626614
rect 372954 590614 373574 626058
rect 372954 590058 372986 590614
rect 373542 590058 373574 590614
rect 372954 554614 373574 590058
rect 372954 554058 372986 554614
rect 373542 554058 373574 554614
rect 372954 518614 373574 554058
rect 372954 518058 372986 518614
rect 373542 518058 373574 518614
rect 372954 482614 373574 518058
rect 372954 482058 372986 482614
rect 373542 482058 373574 482614
rect 372954 460000 373574 482058
rect 379794 705798 380414 705830
rect 379794 705242 379826 705798
rect 380382 705242 380414 705798
rect 379794 669454 380414 705242
rect 379794 668898 379826 669454
rect 380382 668898 380414 669454
rect 379794 633454 380414 668898
rect 379794 632898 379826 633454
rect 380382 632898 380414 633454
rect 379794 597454 380414 632898
rect 379794 596898 379826 597454
rect 380382 596898 380414 597454
rect 379794 561454 380414 596898
rect 379794 560898 379826 561454
rect 380382 560898 380414 561454
rect 379794 525454 380414 560898
rect 379794 524898 379826 525454
rect 380382 524898 380414 525454
rect 379794 489454 380414 524898
rect 379794 488898 379826 489454
rect 380382 488898 380414 489454
rect 379794 458000 380414 488898
rect 383514 673174 384134 707162
rect 383514 672618 383546 673174
rect 384102 672618 384134 673174
rect 383514 637174 384134 672618
rect 383514 636618 383546 637174
rect 384102 636618 384134 637174
rect 383514 601174 384134 636618
rect 383514 600618 383546 601174
rect 384102 600618 384134 601174
rect 383514 565174 384134 600618
rect 383514 564618 383546 565174
rect 384102 564618 384134 565174
rect 383514 529174 384134 564618
rect 383514 528618 383546 529174
rect 384102 528618 384134 529174
rect 383514 493174 384134 528618
rect 383514 492618 383546 493174
rect 384102 492618 384134 493174
rect 383514 460000 384134 492618
rect 387234 676894 387854 709082
rect 387234 676338 387266 676894
rect 387822 676338 387854 676894
rect 387234 640894 387854 676338
rect 387234 640338 387266 640894
rect 387822 640338 387854 640894
rect 387234 604894 387854 640338
rect 387234 604338 387266 604894
rect 387822 604338 387854 604894
rect 387234 568894 387854 604338
rect 387234 568338 387266 568894
rect 387822 568338 387854 568894
rect 387234 532894 387854 568338
rect 387234 532338 387266 532894
rect 387822 532338 387854 532894
rect 387234 496894 387854 532338
rect 387234 496338 387266 496894
rect 387822 496338 387854 496894
rect 387234 460894 387854 496338
rect 387234 460338 387266 460894
rect 387822 460338 387854 460894
rect 387234 460000 387854 460338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710042 408986 710598
rect 409542 710042 409574 710598
rect 405234 708678 405854 709670
rect 405234 708122 405266 708678
rect 405822 708122 405854 708678
rect 401514 706758 402134 707750
rect 401514 706202 401546 706758
rect 402102 706202 402134 706758
rect 390954 680058 390986 680614
rect 391542 680058 391574 680614
rect 390954 644614 391574 680058
rect 390954 644058 390986 644614
rect 391542 644058 391574 644614
rect 390954 608614 391574 644058
rect 390954 608058 390986 608614
rect 391542 608058 391574 608614
rect 390954 572614 391574 608058
rect 390954 572058 390986 572614
rect 391542 572058 391574 572614
rect 390954 536614 391574 572058
rect 390954 536058 390986 536614
rect 391542 536058 391574 536614
rect 390954 500614 391574 536058
rect 390954 500058 390986 500614
rect 391542 500058 391574 500614
rect 390954 464614 391574 500058
rect 390954 464058 390986 464614
rect 391542 464058 391574 464614
rect 390954 460000 391574 464058
rect 397794 704838 398414 705830
rect 397794 704282 397826 704838
rect 398382 704282 398414 704838
rect 397794 687454 398414 704282
rect 397794 686898 397826 687454
rect 398382 686898 398414 687454
rect 397794 651454 398414 686898
rect 397794 650898 397826 651454
rect 398382 650898 398414 651454
rect 397794 615454 398414 650898
rect 397794 614898 397826 615454
rect 398382 614898 398414 615454
rect 397794 579454 398414 614898
rect 397794 578898 397826 579454
rect 398382 578898 398414 579454
rect 397794 543454 398414 578898
rect 397794 542898 397826 543454
rect 398382 542898 398414 543454
rect 397794 507454 398414 542898
rect 397794 506898 397826 507454
rect 398382 506898 398414 507454
rect 397794 471454 398414 506898
rect 397794 470898 397826 471454
rect 398382 470898 398414 471454
rect 397794 458000 398414 470898
rect 401514 691174 402134 706202
rect 401514 690618 401546 691174
rect 402102 690618 402134 691174
rect 401514 655174 402134 690618
rect 401514 654618 401546 655174
rect 402102 654618 402134 655174
rect 401514 619174 402134 654618
rect 401514 618618 401546 619174
rect 402102 618618 402134 619174
rect 401514 583174 402134 618618
rect 401514 582618 401546 583174
rect 402102 582618 402134 583174
rect 401514 547174 402134 582618
rect 401514 546618 401546 547174
rect 402102 546618 402134 547174
rect 401514 511174 402134 546618
rect 401514 510618 401546 511174
rect 402102 510618 402134 511174
rect 401514 475174 402134 510618
rect 401514 474618 401546 475174
rect 402102 474618 402134 475174
rect 401514 460000 402134 474618
rect 405234 694894 405854 708122
rect 405234 694338 405266 694894
rect 405822 694338 405854 694894
rect 405234 658894 405854 694338
rect 405234 658338 405266 658894
rect 405822 658338 405854 658894
rect 405234 622894 405854 658338
rect 405234 622338 405266 622894
rect 405822 622338 405854 622894
rect 405234 586894 405854 622338
rect 405234 586338 405266 586894
rect 405822 586338 405854 586894
rect 405234 550894 405854 586338
rect 405234 550338 405266 550894
rect 405822 550338 405854 550894
rect 405234 514894 405854 550338
rect 405234 514338 405266 514894
rect 405822 514338 405854 514894
rect 405234 478894 405854 514338
rect 405234 478338 405266 478894
rect 405822 478338 405854 478894
rect 405234 460000 405854 478338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711002 426986 711558
rect 427542 711002 427574 711558
rect 423234 709638 423854 709670
rect 423234 709082 423266 709638
rect 423822 709082 423854 709638
rect 419514 707718 420134 707750
rect 419514 707162 419546 707718
rect 420102 707162 420134 707718
rect 408954 698058 408986 698614
rect 409542 698058 409574 698614
rect 408954 662614 409574 698058
rect 408954 662058 408986 662614
rect 409542 662058 409574 662614
rect 408954 626614 409574 662058
rect 408954 626058 408986 626614
rect 409542 626058 409574 626614
rect 408954 590614 409574 626058
rect 408954 590058 408986 590614
rect 409542 590058 409574 590614
rect 408954 554614 409574 590058
rect 408954 554058 408986 554614
rect 409542 554058 409574 554614
rect 408954 518614 409574 554058
rect 408954 518058 408986 518614
rect 409542 518058 409574 518614
rect 408954 482614 409574 518058
rect 408954 482058 408986 482614
rect 409542 482058 409574 482614
rect 408954 460000 409574 482058
rect 415794 705798 416414 705830
rect 415794 705242 415826 705798
rect 416382 705242 416414 705798
rect 415794 669454 416414 705242
rect 415794 668898 415826 669454
rect 416382 668898 416414 669454
rect 415794 633454 416414 668898
rect 415794 632898 415826 633454
rect 416382 632898 416414 633454
rect 415794 597454 416414 632898
rect 415794 596898 415826 597454
rect 416382 596898 416414 597454
rect 415794 561454 416414 596898
rect 415794 560898 415826 561454
rect 416382 560898 416414 561454
rect 415794 525454 416414 560898
rect 415794 524898 415826 525454
rect 416382 524898 416414 525454
rect 415794 489454 416414 524898
rect 415794 488898 415826 489454
rect 416382 488898 416414 489454
rect 237235 457332 237301 457333
rect 237235 457268 237236 457332
rect 237300 457268 237301 457332
rect 237235 457267 237301 457268
rect 241283 457332 241349 457333
rect 241283 457268 241284 457332
rect 241348 457268 241349 457332
rect 241283 457267 241349 457268
rect 242755 457332 242821 457333
rect 242755 457268 242756 457332
rect 242820 457268 242821 457332
rect 242755 457267 242821 457268
rect 244043 457332 244109 457333
rect 244043 457268 244044 457332
rect 244108 457268 244109 457332
rect 244043 457267 244109 457268
rect 245515 457332 245581 457333
rect 245515 457268 245516 457332
rect 245580 457268 245581 457332
rect 245515 457267 245581 457268
rect 246803 457332 246869 457333
rect 246803 457268 246804 457332
rect 246868 457268 246869 457332
rect 246803 457267 246869 457268
rect 248275 457332 248341 457333
rect 248275 457268 248276 457332
rect 248340 457268 248341 457332
rect 248275 457267 248341 457268
rect 251035 457332 251101 457333
rect 251035 457268 251036 457332
rect 251100 457268 251101 457332
rect 251035 457267 251101 457268
rect 252323 457332 252389 457333
rect 252323 457268 252324 457332
rect 252388 457268 252389 457332
rect 252323 457267 252389 457268
rect 253611 457332 253677 457333
rect 253611 457268 253612 457332
rect 253676 457268 253677 457332
rect 253611 457267 253677 457268
rect 256555 457332 256621 457333
rect 256555 457268 256556 457332
rect 256620 457268 256621 457332
rect 256555 457267 256621 457268
rect 257291 457332 257357 457333
rect 257291 457268 257292 457332
rect 257356 457268 257357 457332
rect 257291 457267 257357 457268
rect 259315 457332 259381 457333
rect 259315 457268 259316 457332
rect 259380 457268 259381 457332
rect 259315 457267 259381 457268
rect 262075 457332 262141 457333
rect 262075 457268 262076 457332
rect 262140 457268 262141 457332
rect 262075 457267 262141 457268
rect 263363 457332 263429 457333
rect 263363 457268 263364 457332
rect 263428 457268 263429 457332
rect 263363 457267 263429 457268
rect 264651 457332 264717 457333
rect 264651 457268 264652 457332
rect 264716 457268 264717 457332
rect 264651 457267 264717 457268
rect 266123 457332 266189 457333
rect 266123 457268 266124 457332
rect 266188 457268 266189 457332
rect 266123 457267 266189 457268
rect 267595 457332 267661 457333
rect 267595 457268 267596 457332
rect 267660 457268 267661 457332
rect 267595 457267 267661 457268
rect 268883 457332 268949 457333
rect 268883 457268 268884 457332
rect 268948 457268 268949 457332
rect 268883 457267 268949 457268
rect 382227 457332 382293 457333
rect 382227 457268 382228 457332
rect 382292 457268 382293 457332
rect 382227 457267 382293 457268
rect 384251 457332 384317 457333
rect 384251 457268 384252 457332
rect 384316 457268 384317 457332
rect 384251 457267 384317 457268
rect 384987 457332 385053 457333
rect 384987 457268 384988 457332
rect 385052 457268 385053 457332
rect 384987 457267 385053 457268
rect 386459 457332 386525 457333
rect 386459 457268 386460 457332
rect 386524 457268 386525 457332
rect 386459 457267 386525 457268
rect 387931 457332 387997 457333
rect 387931 457268 387932 457332
rect 387996 457268 387997 457332
rect 387931 457267 387997 457268
rect 389219 457332 389285 457333
rect 389219 457268 389220 457332
rect 389284 457268 389285 457332
rect 389219 457267 389285 457268
rect 393451 457332 393517 457333
rect 393451 457268 393452 457332
rect 393516 457268 393517 457332
rect 393451 457267 393517 457268
rect 394739 457332 394805 457333
rect 394739 457268 394740 457332
rect 394804 457268 394805 457332
rect 394739 457267 394805 457268
rect 396211 457332 396277 457333
rect 396211 457268 396212 457332
rect 396276 457268 396277 457332
rect 396211 457267 396277 457268
rect 397499 457332 397565 457333
rect 397499 457268 397500 457332
rect 397564 457268 397565 457332
rect 397499 457267 397565 457268
rect 398787 457332 398853 457333
rect 398787 457268 398788 457332
rect 398852 457268 398853 457332
rect 398787 457267 398853 457268
rect 400259 457332 400325 457333
rect 400259 457268 400260 457332
rect 400324 457268 400325 457332
rect 400259 457267 400325 457268
rect 403019 457332 403085 457333
rect 403019 457268 403020 457332
rect 403084 457268 403085 457332
rect 403019 457267 403085 457268
rect 404307 457332 404373 457333
rect 404307 457268 404308 457332
rect 404372 457268 404373 457332
rect 404307 457267 404373 457268
rect 405963 457332 406029 457333
rect 405963 457268 405964 457332
rect 406028 457268 406029 457332
rect 405963 457267 406029 457268
rect 408723 457332 408789 457333
rect 408723 457268 408724 457332
rect 408788 457268 408789 457332
rect 408723 457267 408789 457268
rect 409827 457332 409893 457333
rect 409827 457268 409828 457332
rect 409892 457268 409893 457332
rect 409827 457267 409893 457268
rect 411299 457332 411365 457333
rect 411299 457268 411300 457332
rect 411364 457268 411365 457332
rect 411299 457267 411365 457268
rect 228954 446058 228986 446614
rect 229542 446058 229574 446614
rect 228954 410614 229574 446058
rect 228954 410058 228986 410614
rect 229542 410058 229574 410614
rect 228954 374614 229574 410058
rect 228954 374058 228986 374614
rect 229542 374058 229574 374614
rect 228954 338614 229574 374058
rect 228954 338058 228986 338614
rect 229542 338058 229574 338614
rect 228954 302614 229574 338058
rect 228954 302058 228986 302614
rect 229542 302058 229574 302614
rect 228954 266614 229574 302058
rect 228954 266058 228986 266614
rect 229542 266058 229574 266614
rect 228954 230614 229574 266058
rect 228954 230058 228986 230614
rect 229542 230058 229574 230614
rect 228954 194614 229574 230058
rect 228954 194058 228986 194614
rect 229542 194058 229574 194614
rect 228954 158614 229574 194058
rect 228954 158058 228986 158614
rect 229542 158058 229574 158614
rect 228954 122614 229574 158058
rect 228954 122058 228986 122614
rect 229542 122058 229574 122614
rect 228954 86614 229574 122058
rect 228954 86058 228986 86614
rect 229542 86058 229574 86614
rect 228954 50614 229574 86058
rect 228954 50058 228986 50614
rect 229542 50058 229574 50614
rect 228954 14614 229574 50058
rect 228954 14058 228986 14614
rect 229542 14058 229574 14614
rect 210954 -7622 210986 -7066
rect 211542 -7622 211574 -7066
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 309454 236414 338000
rect 235794 308898 235826 309454
rect 236382 308898 236414 309454
rect 235794 273454 236414 308898
rect 235794 272898 235826 273454
rect 236382 272898 236414 273454
rect 235794 237454 236414 272898
rect 235794 236898 235826 237454
rect 236382 236898 236414 237454
rect 235794 201454 236414 236898
rect 235794 200898 235826 201454
rect 236382 200898 236414 201454
rect 235794 165454 236414 200898
rect 235794 164898 235826 165454
rect 236382 164898 236414 165454
rect 235794 129454 236414 164898
rect 235794 128898 235826 129454
rect 236382 128898 236414 129454
rect 235794 93454 236414 128898
rect 235794 92898 235826 93454
rect 236382 92898 236414 93454
rect 235794 57454 236414 92898
rect 235794 56898 235826 57454
rect 236382 56898 236414 57454
rect 235794 21454 236414 56898
rect 237238 31789 237298 457267
rect 239208 435454 239528 435486
rect 239208 435218 239250 435454
rect 239486 435218 239528 435454
rect 239208 435134 239528 435218
rect 239208 434898 239250 435134
rect 239486 434898 239528 435134
rect 239208 434866 239528 434898
rect 239208 399454 239528 399486
rect 239208 399218 239250 399454
rect 239486 399218 239528 399454
rect 239208 399134 239528 399218
rect 239208 398898 239250 399134
rect 239486 398898 239528 399134
rect 239208 398866 239528 398898
rect 239208 363454 239528 363486
rect 239208 363218 239250 363454
rect 239486 363218 239528 363454
rect 239208 363134 239528 363218
rect 239208 362898 239250 363134
rect 239486 362898 239528 363134
rect 239208 362866 239528 362898
rect 239514 313174 240134 336000
rect 239514 312618 239546 313174
rect 240102 312618 240134 313174
rect 239514 277174 240134 312618
rect 239514 276618 239546 277174
rect 240102 276618 240134 277174
rect 239514 241174 240134 276618
rect 239514 240618 239546 241174
rect 240102 240618 240134 241174
rect 239514 205174 240134 240618
rect 239514 204618 239546 205174
rect 240102 204618 240134 205174
rect 239514 169174 240134 204618
rect 239514 168618 239546 169174
rect 240102 168618 240134 169174
rect 239514 133174 240134 168618
rect 239514 132618 239546 133174
rect 240102 132618 240134 133174
rect 239514 97174 240134 132618
rect 239514 96618 239546 97174
rect 240102 96618 240134 97174
rect 239514 61174 240134 96618
rect 239514 60618 239546 61174
rect 240102 60618 240134 61174
rect 237235 31788 237301 31789
rect 237235 31724 237236 31788
rect 237300 31724 237301 31788
rect 237235 31723 237301 31724
rect 235794 20898 235826 21454
rect 236382 20898 236414 21454
rect 235794 -1306 236414 20898
rect 235794 -1862 235826 -1306
rect 236382 -1862 236414 -1306
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 60618
rect 241286 45661 241346 457267
rect 242758 71909 242818 457267
rect 243234 316894 243854 336000
rect 243234 316338 243266 316894
rect 243822 316338 243854 316894
rect 243234 280894 243854 316338
rect 243234 280338 243266 280894
rect 243822 280338 243854 280894
rect 243234 244894 243854 280338
rect 243234 244338 243266 244894
rect 243822 244338 243854 244894
rect 243234 208894 243854 244338
rect 243234 208338 243266 208894
rect 243822 208338 243854 208894
rect 243234 172894 243854 208338
rect 243234 172338 243266 172894
rect 243822 172338 243854 172894
rect 243234 136894 243854 172338
rect 243234 136338 243266 136894
rect 243822 136338 243854 136894
rect 243234 100894 243854 136338
rect 243234 100338 243266 100894
rect 243822 100338 243854 100894
rect 242755 71908 242821 71909
rect 242755 71844 242756 71908
rect 242820 71844 242821 71908
rect 242755 71843 242821 71844
rect 243234 64894 243854 100338
rect 243234 64338 243266 64894
rect 243822 64338 243854 64894
rect 241283 45660 241349 45661
rect 241283 45596 241284 45660
rect 241348 45596 241349 45660
rect 241283 45595 241349 45596
rect 239514 24618 239546 25174
rect 240102 24618 240134 25174
rect 239514 -3226 240134 24618
rect 239514 -3782 239546 -3226
rect 240102 -3782 240134 -3226
rect 239514 -3814 240134 -3782
rect 243234 28894 243854 64338
rect 244046 59397 244106 457267
rect 245518 85645 245578 457267
rect 246806 111893 246866 457267
rect 246954 320614 247574 336000
rect 246954 320058 246986 320614
rect 247542 320058 247574 320614
rect 246954 284614 247574 320058
rect 246954 284058 246986 284614
rect 247542 284058 247574 284614
rect 246954 248614 247574 284058
rect 246954 248058 246986 248614
rect 247542 248058 247574 248614
rect 246954 212614 247574 248058
rect 246954 212058 246986 212614
rect 247542 212058 247574 212614
rect 246954 176614 247574 212058
rect 246954 176058 246986 176614
rect 247542 176058 247574 176614
rect 246954 140614 247574 176058
rect 246954 140058 246986 140614
rect 247542 140058 247574 140614
rect 246803 111892 246869 111893
rect 246803 111828 246804 111892
rect 246868 111828 246869 111892
rect 246803 111827 246869 111828
rect 246954 104614 247574 140058
rect 246954 104058 246986 104614
rect 247542 104058 247574 104614
rect 245515 85644 245581 85645
rect 245515 85580 245516 85644
rect 245580 85580 245581 85644
rect 245515 85579 245581 85580
rect 246954 68614 247574 104058
rect 248278 99517 248338 457267
rect 251038 125629 251098 457267
rect 252326 151877 252386 457267
rect 252323 151876 252389 151877
rect 252323 151812 252324 151876
rect 252388 151812 252389 151876
rect 252323 151811 252389 151812
rect 253614 138141 253674 457267
rect 254568 453454 254888 453486
rect 254568 453218 254610 453454
rect 254846 453218 254888 453454
rect 254568 453134 254888 453218
rect 254568 452898 254610 453134
rect 254846 452898 254888 453134
rect 254568 452866 254888 452898
rect 254568 417454 254888 417486
rect 254568 417218 254610 417454
rect 254846 417218 254888 417454
rect 254568 417134 254888 417218
rect 254568 416898 254610 417134
rect 254846 416898 254888 417134
rect 254568 416866 254888 416898
rect 254568 381454 254888 381486
rect 254568 381218 254610 381454
rect 254846 381218 254888 381454
rect 254568 381134 254888 381218
rect 254568 380898 254610 381134
rect 254846 380898 254888 381134
rect 254568 380866 254888 380898
rect 254568 345454 254888 345486
rect 254568 345218 254610 345454
rect 254846 345218 254888 345454
rect 254568 345134 254888 345218
rect 254568 344898 254610 345134
rect 254846 344898 254888 345134
rect 254568 344866 254888 344898
rect 253794 327454 254414 338000
rect 253794 326898 253826 327454
rect 254382 326898 254414 327454
rect 253794 291454 254414 326898
rect 253794 290898 253826 291454
rect 254382 290898 254414 291454
rect 253794 255454 254414 290898
rect 253794 254898 253826 255454
rect 254382 254898 254414 255454
rect 253794 219454 254414 254898
rect 253794 218898 253826 219454
rect 254382 218898 254414 219454
rect 253794 183454 254414 218898
rect 256558 191861 256618 457267
rect 256555 191860 256621 191861
rect 256555 191796 256556 191860
rect 256620 191796 256621 191860
rect 256555 191795 256621 191796
rect 253794 182898 253826 183454
rect 254382 182898 254414 183454
rect 253794 147454 254414 182898
rect 257294 178125 257354 457267
rect 257514 331174 258134 336000
rect 257514 330618 257546 331174
rect 258102 330618 258134 331174
rect 257514 295174 258134 330618
rect 257514 294618 257546 295174
rect 258102 294618 258134 295174
rect 257514 259174 258134 294618
rect 257514 258618 257546 259174
rect 258102 258618 258134 259174
rect 257514 223174 258134 258618
rect 257514 222618 257546 223174
rect 258102 222618 258134 223174
rect 257514 187174 258134 222618
rect 259318 205733 259378 457267
rect 261234 334894 261854 336000
rect 261234 334338 261266 334894
rect 261822 334338 261854 334894
rect 261234 298894 261854 334338
rect 261234 298338 261266 298894
rect 261822 298338 261854 298894
rect 261234 262894 261854 298338
rect 261234 262338 261266 262894
rect 261822 262338 261854 262894
rect 261234 226894 261854 262338
rect 262078 231981 262138 457267
rect 262075 231980 262141 231981
rect 262075 231916 262076 231980
rect 262140 231916 262141 231980
rect 262075 231915 262141 231916
rect 261234 226338 261266 226894
rect 261822 226338 261854 226894
rect 259315 205732 259381 205733
rect 259315 205668 259316 205732
rect 259380 205668 259381 205732
rect 259315 205667 259381 205668
rect 257514 186618 257546 187174
rect 258102 186618 258134 187174
rect 257291 178124 257357 178125
rect 257291 178060 257292 178124
rect 257356 178060 257357 178124
rect 257291 178059 257357 178060
rect 253794 146898 253826 147454
rect 254382 146898 254414 147454
rect 253611 138140 253677 138141
rect 253611 138076 253612 138140
rect 253676 138076 253677 138140
rect 253611 138075 253677 138076
rect 251035 125628 251101 125629
rect 251035 125564 251036 125628
rect 251100 125564 251101 125628
rect 251035 125563 251101 125564
rect 253794 111454 254414 146898
rect 253794 110898 253826 111454
rect 254382 110898 254414 111454
rect 248275 99516 248341 99517
rect 248275 99452 248276 99516
rect 248340 99452 248341 99516
rect 248275 99451 248341 99452
rect 246954 68058 246986 68614
rect 247542 68058 247574 68614
rect 244043 59396 244109 59397
rect 244043 59332 244044 59396
rect 244108 59332 244109 59396
rect 244043 59331 244109 59332
rect 243234 28338 243266 28894
rect 243822 28338 243854 28894
rect 243234 -5146 243854 28338
rect 243234 -5702 243266 -5146
rect 243822 -5702 243854 -5146
rect 243234 -5734 243854 -5702
rect 246954 32614 247574 68058
rect 246954 32058 246986 32614
rect 247542 32058 247574 32614
rect 228954 -6662 228986 -6106
rect 229542 -6662 229574 -6106
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 75454 254414 110898
rect 253794 74898 253826 75454
rect 254382 74898 254414 75454
rect 253794 39454 254414 74898
rect 253794 38898 253826 39454
rect 254382 38898 254414 39454
rect 253794 3454 254414 38898
rect 253794 2898 253826 3454
rect 254382 2898 254414 3454
rect 253794 -346 254414 2898
rect 253794 -902 253826 -346
rect 254382 -902 254414 -346
rect 253794 -1894 254414 -902
rect 257514 151174 258134 186618
rect 257514 150618 257546 151174
rect 258102 150618 258134 151174
rect 257514 115174 258134 150618
rect 257514 114618 257546 115174
rect 258102 114618 258134 115174
rect 257514 79174 258134 114618
rect 257514 78618 257546 79174
rect 258102 78618 258134 79174
rect 257514 43174 258134 78618
rect 257514 42618 257546 43174
rect 258102 42618 258134 43174
rect 257514 7174 258134 42618
rect 257514 6618 257546 7174
rect 258102 6618 258134 7174
rect 257514 -2266 258134 6618
rect 257514 -2822 257546 -2266
rect 258102 -2822 258134 -2266
rect 257514 -3814 258134 -2822
rect 261234 190894 261854 226338
rect 263366 218109 263426 457267
rect 264654 244357 264714 457267
rect 264954 302614 265574 336000
rect 264954 302058 264986 302614
rect 265542 302058 265574 302614
rect 264954 266614 265574 302058
rect 266126 271965 266186 457267
rect 266123 271964 266189 271965
rect 266123 271900 266124 271964
rect 266188 271900 266189 271964
rect 266123 271899 266189 271900
rect 264954 266058 264986 266614
rect 265542 266058 265574 266614
rect 264651 244356 264717 244357
rect 264651 244292 264652 244356
rect 264716 244292 264717 244356
rect 264651 244291 264717 244292
rect 264954 230614 265574 266058
rect 267598 258093 267658 457267
rect 268886 298213 268946 457267
rect 285288 453454 285608 453486
rect 285288 453218 285330 453454
rect 285566 453218 285608 453454
rect 285288 453134 285608 453218
rect 285288 452898 285330 453134
rect 285566 452898 285608 453134
rect 285288 452866 285608 452898
rect 316008 453454 316328 453486
rect 316008 453218 316050 453454
rect 316286 453218 316328 453454
rect 316008 453134 316328 453218
rect 316008 452898 316050 453134
rect 316286 452898 316328 453134
rect 316008 452866 316328 452898
rect 346728 453454 347048 453486
rect 346728 453218 346770 453454
rect 347006 453218 347048 453454
rect 346728 453134 347048 453218
rect 346728 452898 346770 453134
rect 347006 452898 347048 453134
rect 346728 452866 347048 452898
rect 377448 453454 377768 453486
rect 377448 453218 377490 453454
rect 377726 453218 377768 453454
rect 377448 453134 377768 453218
rect 377448 452898 377490 453134
rect 377726 452898 377768 453134
rect 377448 452866 377768 452898
rect 269928 435454 270248 435486
rect 269928 435218 269970 435454
rect 270206 435218 270248 435454
rect 269928 435134 270248 435218
rect 269928 434898 269970 435134
rect 270206 434898 270248 435134
rect 269928 434866 270248 434898
rect 300648 435454 300968 435486
rect 300648 435218 300690 435454
rect 300926 435218 300968 435454
rect 300648 435134 300968 435218
rect 300648 434898 300690 435134
rect 300926 434898 300968 435134
rect 300648 434866 300968 434898
rect 331368 435454 331688 435486
rect 331368 435218 331410 435454
rect 331646 435218 331688 435454
rect 331368 435134 331688 435218
rect 331368 434898 331410 435134
rect 331646 434898 331688 435134
rect 331368 434866 331688 434898
rect 362088 435454 362408 435486
rect 362088 435218 362130 435454
rect 362366 435218 362408 435454
rect 362088 435134 362408 435218
rect 362088 434898 362130 435134
rect 362366 434898 362408 435134
rect 362088 434866 362408 434898
rect 285288 417454 285608 417486
rect 285288 417218 285330 417454
rect 285566 417218 285608 417454
rect 285288 417134 285608 417218
rect 285288 416898 285330 417134
rect 285566 416898 285608 417134
rect 285288 416866 285608 416898
rect 316008 417454 316328 417486
rect 316008 417218 316050 417454
rect 316286 417218 316328 417454
rect 316008 417134 316328 417218
rect 316008 416898 316050 417134
rect 316286 416898 316328 417134
rect 316008 416866 316328 416898
rect 346728 417454 347048 417486
rect 346728 417218 346770 417454
rect 347006 417218 347048 417454
rect 346728 417134 347048 417218
rect 346728 416898 346770 417134
rect 347006 416898 347048 417134
rect 346728 416866 347048 416898
rect 377448 417454 377768 417486
rect 377448 417218 377490 417454
rect 377726 417218 377768 417454
rect 377448 417134 377768 417218
rect 377448 416898 377490 417134
rect 377726 416898 377768 417134
rect 377448 416866 377768 416898
rect 269928 399454 270248 399486
rect 269928 399218 269970 399454
rect 270206 399218 270248 399454
rect 269928 399134 270248 399218
rect 269928 398898 269970 399134
rect 270206 398898 270248 399134
rect 269928 398866 270248 398898
rect 300648 399454 300968 399486
rect 300648 399218 300690 399454
rect 300926 399218 300968 399454
rect 300648 399134 300968 399218
rect 300648 398898 300690 399134
rect 300926 398898 300968 399134
rect 300648 398866 300968 398898
rect 331368 399454 331688 399486
rect 331368 399218 331410 399454
rect 331646 399218 331688 399454
rect 331368 399134 331688 399218
rect 331368 398898 331410 399134
rect 331646 398898 331688 399134
rect 331368 398866 331688 398898
rect 362088 399454 362408 399486
rect 362088 399218 362130 399454
rect 362366 399218 362408 399454
rect 362088 399134 362408 399218
rect 362088 398898 362130 399134
rect 362366 398898 362408 399134
rect 362088 398866 362408 398898
rect 285288 381454 285608 381486
rect 285288 381218 285330 381454
rect 285566 381218 285608 381454
rect 285288 381134 285608 381218
rect 285288 380898 285330 381134
rect 285566 380898 285608 381134
rect 285288 380866 285608 380898
rect 316008 381454 316328 381486
rect 316008 381218 316050 381454
rect 316286 381218 316328 381454
rect 316008 381134 316328 381218
rect 316008 380898 316050 381134
rect 316286 380898 316328 381134
rect 316008 380866 316328 380898
rect 346728 381454 347048 381486
rect 346728 381218 346770 381454
rect 347006 381218 347048 381454
rect 346728 381134 347048 381218
rect 346728 380898 346770 381134
rect 347006 380898 347048 381134
rect 346728 380866 347048 380898
rect 377448 381454 377768 381486
rect 377448 381218 377490 381454
rect 377726 381218 377768 381454
rect 377448 381134 377768 381218
rect 377448 380898 377490 381134
rect 377726 380898 377768 381134
rect 377448 380866 377768 380898
rect 269928 363454 270248 363486
rect 269928 363218 269970 363454
rect 270206 363218 270248 363454
rect 269928 363134 270248 363218
rect 269928 362898 269970 363134
rect 270206 362898 270248 363134
rect 269928 362866 270248 362898
rect 300648 363454 300968 363486
rect 300648 363218 300690 363454
rect 300926 363218 300968 363454
rect 300648 363134 300968 363218
rect 300648 362898 300690 363134
rect 300926 362898 300968 363134
rect 300648 362866 300968 362898
rect 331368 363454 331688 363486
rect 331368 363218 331410 363454
rect 331646 363218 331688 363454
rect 331368 363134 331688 363218
rect 331368 362898 331410 363134
rect 331646 362898 331688 363134
rect 331368 362866 331688 362898
rect 362088 363454 362408 363486
rect 362088 363218 362130 363454
rect 362366 363218 362408 363454
rect 362088 363134 362408 363218
rect 362088 362898 362130 363134
rect 362366 362898 362408 363134
rect 362088 362866 362408 362898
rect 285288 345454 285608 345486
rect 285288 345218 285330 345454
rect 285566 345218 285608 345454
rect 285288 345134 285608 345218
rect 285288 344898 285330 345134
rect 285566 344898 285608 345134
rect 285288 344866 285608 344898
rect 316008 345454 316328 345486
rect 316008 345218 316050 345454
rect 316286 345218 316328 345454
rect 316008 345134 316328 345218
rect 316008 344898 316050 345134
rect 316286 344898 316328 345134
rect 316008 344866 316328 344898
rect 346728 345454 347048 345486
rect 346728 345218 346770 345454
rect 347006 345218 347048 345454
rect 346728 345134 347048 345218
rect 346728 344898 346770 345134
rect 347006 344898 347048 345134
rect 346728 344866 347048 344898
rect 377448 345454 377768 345486
rect 377448 345218 377490 345454
rect 377726 345218 377768 345454
rect 377448 345134 377768 345218
rect 377448 344898 377490 345134
rect 377726 344898 377768 345134
rect 377448 344866 377768 344898
rect 271794 309454 272414 338000
rect 271794 308898 271826 309454
rect 272382 308898 272414 309454
rect 268883 298212 268949 298213
rect 268883 298148 268884 298212
rect 268948 298148 268949 298212
rect 268883 298147 268949 298148
rect 271794 273454 272414 308898
rect 271794 272898 271826 273454
rect 272382 272898 272414 273454
rect 267595 258092 267661 258093
rect 267595 258028 267596 258092
rect 267660 258028 267661 258092
rect 267595 258027 267661 258028
rect 264954 230058 264986 230614
rect 265542 230058 265574 230614
rect 263363 218108 263429 218109
rect 263363 218044 263364 218108
rect 263428 218044 263429 218108
rect 263363 218043 263429 218044
rect 261234 190338 261266 190894
rect 261822 190338 261854 190894
rect 261234 154894 261854 190338
rect 261234 154338 261266 154894
rect 261822 154338 261854 154894
rect 261234 118894 261854 154338
rect 261234 118338 261266 118894
rect 261822 118338 261854 118894
rect 261234 82894 261854 118338
rect 261234 82338 261266 82894
rect 261822 82338 261854 82894
rect 261234 46894 261854 82338
rect 261234 46338 261266 46894
rect 261822 46338 261854 46894
rect 261234 10894 261854 46338
rect 261234 10338 261266 10894
rect 261822 10338 261854 10894
rect 261234 -4186 261854 10338
rect 261234 -4742 261266 -4186
rect 261822 -4742 261854 -4186
rect 261234 -5734 261854 -4742
rect 264954 194614 265574 230058
rect 264954 194058 264986 194614
rect 265542 194058 265574 194614
rect 264954 158614 265574 194058
rect 264954 158058 264986 158614
rect 265542 158058 265574 158614
rect 264954 122614 265574 158058
rect 264954 122058 264986 122614
rect 265542 122058 265574 122614
rect 264954 86614 265574 122058
rect 264954 86058 264986 86614
rect 265542 86058 265574 86614
rect 264954 50614 265574 86058
rect 264954 50058 264986 50614
rect 265542 50058 265574 50614
rect 264954 14614 265574 50058
rect 264954 14058 264986 14614
rect 265542 14058 265574 14614
rect 246954 -7622 246986 -7066
rect 247542 -7622 247574 -7066
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 237454 272414 272898
rect 271794 236898 271826 237454
rect 272382 236898 272414 237454
rect 271794 201454 272414 236898
rect 271794 200898 271826 201454
rect 272382 200898 272414 201454
rect 271794 165454 272414 200898
rect 271794 164898 271826 165454
rect 272382 164898 272414 165454
rect 271794 129454 272414 164898
rect 271794 128898 271826 129454
rect 272382 128898 272414 129454
rect 271794 93454 272414 128898
rect 271794 92898 271826 93454
rect 272382 92898 272414 93454
rect 271794 57454 272414 92898
rect 271794 56898 271826 57454
rect 272382 56898 272414 57454
rect 271794 21454 272414 56898
rect 271794 20898 271826 21454
rect 272382 20898 272414 21454
rect 271794 -1306 272414 20898
rect 271794 -1862 271826 -1306
rect 272382 -1862 272414 -1306
rect 271794 -1894 272414 -1862
rect 275514 313174 276134 336000
rect 275514 312618 275546 313174
rect 276102 312618 276134 313174
rect 275514 277174 276134 312618
rect 275514 276618 275546 277174
rect 276102 276618 276134 277174
rect 275514 241174 276134 276618
rect 275514 240618 275546 241174
rect 276102 240618 276134 241174
rect 275514 205174 276134 240618
rect 275514 204618 275546 205174
rect 276102 204618 276134 205174
rect 275514 169174 276134 204618
rect 275514 168618 275546 169174
rect 276102 168618 276134 169174
rect 275514 133174 276134 168618
rect 275514 132618 275546 133174
rect 276102 132618 276134 133174
rect 275514 97174 276134 132618
rect 275514 96618 275546 97174
rect 276102 96618 276134 97174
rect 275514 61174 276134 96618
rect 275514 60618 275546 61174
rect 276102 60618 276134 61174
rect 275514 25174 276134 60618
rect 275514 24618 275546 25174
rect 276102 24618 276134 25174
rect 275514 -3226 276134 24618
rect 275514 -3782 275546 -3226
rect 276102 -3782 276134 -3226
rect 275514 -3814 276134 -3782
rect 279234 316894 279854 336000
rect 279234 316338 279266 316894
rect 279822 316338 279854 316894
rect 279234 280894 279854 316338
rect 279234 280338 279266 280894
rect 279822 280338 279854 280894
rect 279234 244894 279854 280338
rect 279234 244338 279266 244894
rect 279822 244338 279854 244894
rect 279234 208894 279854 244338
rect 279234 208338 279266 208894
rect 279822 208338 279854 208894
rect 279234 172894 279854 208338
rect 279234 172338 279266 172894
rect 279822 172338 279854 172894
rect 279234 136894 279854 172338
rect 279234 136338 279266 136894
rect 279822 136338 279854 136894
rect 279234 100894 279854 136338
rect 279234 100338 279266 100894
rect 279822 100338 279854 100894
rect 279234 64894 279854 100338
rect 279234 64338 279266 64894
rect 279822 64338 279854 64894
rect 279234 28894 279854 64338
rect 279234 28338 279266 28894
rect 279822 28338 279854 28894
rect 279234 -5146 279854 28338
rect 279234 -5702 279266 -5146
rect 279822 -5702 279854 -5146
rect 279234 -5734 279854 -5702
rect 282954 320614 283574 336000
rect 282954 320058 282986 320614
rect 283542 320058 283574 320614
rect 282954 284614 283574 320058
rect 282954 284058 282986 284614
rect 283542 284058 283574 284614
rect 282954 248614 283574 284058
rect 282954 248058 282986 248614
rect 283542 248058 283574 248614
rect 282954 212614 283574 248058
rect 282954 212058 282986 212614
rect 283542 212058 283574 212614
rect 282954 176614 283574 212058
rect 282954 176058 282986 176614
rect 283542 176058 283574 176614
rect 282954 140614 283574 176058
rect 282954 140058 282986 140614
rect 283542 140058 283574 140614
rect 282954 104614 283574 140058
rect 282954 104058 282986 104614
rect 283542 104058 283574 104614
rect 282954 68614 283574 104058
rect 282954 68058 282986 68614
rect 283542 68058 283574 68614
rect 282954 32614 283574 68058
rect 282954 32058 282986 32614
rect 283542 32058 283574 32614
rect 264954 -6662 264986 -6106
rect 265542 -6662 265574 -6106
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 327454 290414 338000
rect 289794 326898 289826 327454
rect 290382 326898 290414 327454
rect 289794 291454 290414 326898
rect 289794 290898 289826 291454
rect 290382 290898 290414 291454
rect 289794 255454 290414 290898
rect 289794 254898 289826 255454
rect 290382 254898 290414 255454
rect 289794 219454 290414 254898
rect 289794 218898 289826 219454
rect 290382 218898 290414 219454
rect 289794 183454 290414 218898
rect 289794 182898 289826 183454
rect 290382 182898 290414 183454
rect 289794 147454 290414 182898
rect 289794 146898 289826 147454
rect 290382 146898 290414 147454
rect 289794 111454 290414 146898
rect 289794 110898 289826 111454
rect 290382 110898 290414 111454
rect 289794 75454 290414 110898
rect 289794 74898 289826 75454
rect 290382 74898 290414 75454
rect 289794 39454 290414 74898
rect 289794 38898 289826 39454
rect 290382 38898 290414 39454
rect 289794 3454 290414 38898
rect 289794 2898 289826 3454
rect 290382 2898 290414 3454
rect 289794 -346 290414 2898
rect 289794 -902 289826 -346
rect 290382 -902 290414 -346
rect 289794 -1894 290414 -902
rect 293514 331174 294134 336000
rect 293514 330618 293546 331174
rect 294102 330618 294134 331174
rect 293514 295174 294134 330618
rect 293514 294618 293546 295174
rect 294102 294618 294134 295174
rect 293514 259174 294134 294618
rect 293514 258618 293546 259174
rect 294102 258618 294134 259174
rect 293514 223174 294134 258618
rect 293514 222618 293546 223174
rect 294102 222618 294134 223174
rect 293514 187174 294134 222618
rect 293514 186618 293546 187174
rect 294102 186618 294134 187174
rect 293514 151174 294134 186618
rect 293514 150618 293546 151174
rect 294102 150618 294134 151174
rect 293514 115174 294134 150618
rect 293514 114618 293546 115174
rect 294102 114618 294134 115174
rect 293514 79174 294134 114618
rect 293514 78618 293546 79174
rect 294102 78618 294134 79174
rect 293514 43174 294134 78618
rect 293514 42618 293546 43174
rect 294102 42618 294134 43174
rect 293514 7174 294134 42618
rect 293514 6618 293546 7174
rect 294102 6618 294134 7174
rect 293514 -2266 294134 6618
rect 293514 -2822 293546 -2266
rect 294102 -2822 294134 -2266
rect 293514 -3814 294134 -2822
rect 297234 334894 297854 336000
rect 297234 334338 297266 334894
rect 297822 334338 297854 334894
rect 297234 298894 297854 334338
rect 297234 298338 297266 298894
rect 297822 298338 297854 298894
rect 297234 262894 297854 298338
rect 297234 262338 297266 262894
rect 297822 262338 297854 262894
rect 297234 226894 297854 262338
rect 297234 226338 297266 226894
rect 297822 226338 297854 226894
rect 297234 190894 297854 226338
rect 297234 190338 297266 190894
rect 297822 190338 297854 190894
rect 297234 154894 297854 190338
rect 297234 154338 297266 154894
rect 297822 154338 297854 154894
rect 297234 118894 297854 154338
rect 297234 118338 297266 118894
rect 297822 118338 297854 118894
rect 297234 82894 297854 118338
rect 297234 82338 297266 82894
rect 297822 82338 297854 82894
rect 297234 46894 297854 82338
rect 297234 46338 297266 46894
rect 297822 46338 297854 46894
rect 297234 10894 297854 46338
rect 297234 10338 297266 10894
rect 297822 10338 297854 10894
rect 297234 -4186 297854 10338
rect 297234 -4742 297266 -4186
rect 297822 -4742 297854 -4186
rect 297234 -5734 297854 -4742
rect 300954 302614 301574 336000
rect 300954 302058 300986 302614
rect 301542 302058 301574 302614
rect 300954 266614 301574 302058
rect 300954 266058 300986 266614
rect 301542 266058 301574 266614
rect 300954 230614 301574 266058
rect 300954 230058 300986 230614
rect 301542 230058 301574 230614
rect 300954 194614 301574 230058
rect 300954 194058 300986 194614
rect 301542 194058 301574 194614
rect 300954 158614 301574 194058
rect 300954 158058 300986 158614
rect 301542 158058 301574 158614
rect 300954 122614 301574 158058
rect 300954 122058 300986 122614
rect 301542 122058 301574 122614
rect 300954 86614 301574 122058
rect 300954 86058 300986 86614
rect 301542 86058 301574 86614
rect 300954 50614 301574 86058
rect 300954 50058 300986 50614
rect 301542 50058 301574 50614
rect 300954 14614 301574 50058
rect 300954 14058 300986 14614
rect 301542 14058 301574 14614
rect 282954 -7622 282986 -7066
rect 283542 -7622 283574 -7066
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 309454 308414 338000
rect 307794 308898 307826 309454
rect 308382 308898 308414 309454
rect 307794 273454 308414 308898
rect 307794 272898 307826 273454
rect 308382 272898 308414 273454
rect 307794 237454 308414 272898
rect 307794 236898 307826 237454
rect 308382 236898 308414 237454
rect 307794 201454 308414 236898
rect 307794 200898 307826 201454
rect 308382 200898 308414 201454
rect 307794 165454 308414 200898
rect 307794 164898 307826 165454
rect 308382 164898 308414 165454
rect 307794 129454 308414 164898
rect 307794 128898 307826 129454
rect 308382 128898 308414 129454
rect 307794 93454 308414 128898
rect 307794 92898 307826 93454
rect 308382 92898 308414 93454
rect 307794 57454 308414 92898
rect 307794 56898 307826 57454
rect 308382 56898 308414 57454
rect 307794 21454 308414 56898
rect 307794 20898 307826 21454
rect 308382 20898 308414 21454
rect 307794 -1306 308414 20898
rect 307794 -1862 307826 -1306
rect 308382 -1862 308414 -1306
rect 307794 -1894 308414 -1862
rect 311514 313174 312134 336000
rect 311514 312618 311546 313174
rect 312102 312618 312134 313174
rect 311514 277174 312134 312618
rect 311514 276618 311546 277174
rect 312102 276618 312134 277174
rect 311514 241174 312134 276618
rect 311514 240618 311546 241174
rect 312102 240618 312134 241174
rect 311514 205174 312134 240618
rect 311514 204618 311546 205174
rect 312102 204618 312134 205174
rect 311514 169174 312134 204618
rect 311514 168618 311546 169174
rect 312102 168618 312134 169174
rect 311514 133174 312134 168618
rect 311514 132618 311546 133174
rect 312102 132618 312134 133174
rect 311514 97174 312134 132618
rect 311514 96618 311546 97174
rect 312102 96618 312134 97174
rect 311514 61174 312134 96618
rect 311514 60618 311546 61174
rect 312102 60618 312134 61174
rect 311514 25174 312134 60618
rect 311514 24618 311546 25174
rect 312102 24618 312134 25174
rect 311514 -3226 312134 24618
rect 311514 -3782 311546 -3226
rect 312102 -3782 312134 -3226
rect 311514 -3814 312134 -3782
rect 315234 316894 315854 336000
rect 315234 316338 315266 316894
rect 315822 316338 315854 316894
rect 315234 280894 315854 316338
rect 315234 280338 315266 280894
rect 315822 280338 315854 280894
rect 315234 244894 315854 280338
rect 315234 244338 315266 244894
rect 315822 244338 315854 244894
rect 315234 208894 315854 244338
rect 315234 208338 315266 208894
rect 315822 208338 315854 208894
rect 315234 172894 315854 208338
rect 315234 172338 315266 172894
rect 315822 172338 315854 172894
rect 315234 136894 315854 172338
rect 315234 136338 315266 136894
rect 315822 136338 315854 136894
rect 315234 100894 315854 136338
rect 315234 100338 315266 100894
rect 315822 100338 315854 100894
rect 315234 64894 315854 100338
rect 315234 64338 315266 64894
rect 315822 64338 315854 64894
rect 315234 28894 315854 64338
rect 315234 28338 315266 28894
rect 315822 28338 315854 28894
rect 315234 -5146 315854 28338
rect 315234 -5702 315266 -5146
rect 315822 -5702 315854 -5146
rect 315234 -5734 315854 -5702
rect 318954 320614 319574 336000
rect 318954 320058 318986 320614
rect 319542 320058 319574 320614
rect 318954 284614 319574 320058
rect 318954 284058 318986 284614
rect 319542 284058 319574 284614
rect 318954 248614 319574 284058
rect 318954 248058 318986 248614
rect 319542 248058 319574 248614
rect 318954 212614 319574 248058
rect 318954 212058 318986 212614
rect 319542 212058 319574 212614
rect 318954 176614 319574 212058
rect 318954 176058 318986 176614
rect 319542 176058 319574 176614
rect 318954 140614 319574 176058
rect 318954 140058 318986 140614
rect 319542 140058 319574 140614
rect 318954 104614 319574 140058
rect 318954 104058 318986 104614
rect 319542 104058 319574 104614
rect 318954 68614 319574 104058
rect 318954 68058 318986 68614
rect 319542 68058 319574 68614
rect 318954 32614 319574 68058
rect 318954 32058 318986 32614
rect 319542 32058 319574 32614
rect 300954 -6662 300986 -6106
rect 301542 -6662 301574 -6106
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 327454 326414 338000
rect 325794 326898 325826 327454
rect 326382 326898 326414 327454
rect 325794 291454 326414 326898
rect 325794 290898 325826 291454
rect 326382 290898 326414 291454
rect 325794 255454 326414 290898
rect 325794 254898 325826 255454
rect 326382 254898 326414 255454
rect 325794 219454 326414 254898
rect 325794 218898 325826 219454
rect 326382 218898 326414 219454
rect 325794 183454 326414 218898
rect 325794 182898 325826 183454
rect 326382 182898 326414 183454
rect 325794 147454 326414 182898
rect 325794 146898 325826 147454
rect 326382 146898 326414 147454
rect 325794 111454 326414 146898
rect 325794 110898 325826 111454
rect 326382 110898 326414 111454
rect 325794 75454 326414 110898
rect 325794 74898 325826 75454
rect 326382 74898 326414 75454
rect 325794 39454 326414 74898
rect 325794 38898 325826 39454
rect 326382 38898 326414 39454
rect 325794 3454 326414 38898
rect 325794 2898 325826 3454
rect 326382 2898 326414 3454
rect 325794 -346 326414 2898
rect 325794 -902 325826 -346
rect 326382 -902 326414 -346
rect 325794 -1894 326414 -902
rect 329514 331174 330134 336000
rect 329514 330618 329546 331174
rect 330102 330618 330134 331174
rect 329514 295174 330134 330618
rect 329514 294618 329546 295174
rect 330102 294618 330134 295174
rect 329514 259174 330134 294618
rect 329514 258618 329546 259174
rect 330102 258618 330134 259174
rect 329514 223174 330134 258618
rect 329514 222618 329546 223174
rect 330102 222618 330134 223174
rect 329514 187174 330134 222618
rect 329514 186618 329546 187174
rect 330102 186618 330134 187174
rect 329514 151174 330134 186618
rect 329514 150618 329546 151174
rect 330102 150618 330134 151174
rect 329514 115174 330134 150618
rect 329514 114618 329546 115174
rect 330102 114618 330134 115174
rect 329514 79174 330134 114618
rect 329514 78618 329546 79174
rect 330102 78618 330134 79174
rect 329514 43174 330134 78618
rect 329514 42618 329546 43174
rect 330102 42618 330134 43174
rect 329514 7174 330134 42618
rect 329514 6618 329546 7174
rect 330102 6618 330134 7174
rect 329514 -2266 330134 6618
rect 329514 -2822 329546 -2266
rect 330102 -2822 330134 -2266
rect 329514 -3814 330134 -2822
rect 333234 334894 333854 336000
rect 333234 334338 333266 334894
rect 333822 334338 333854 334894
rect 333234 298894 333854 334338
rect 333234 298338 333266 298894
rect 333822 298338 333854 298894
rect 333234 262894 333854 298338
rect 333234 262338 333266 262894
rect 333822 262338 333854 262894
rect 333234 226894 333854 262338
rect 333234 226338 333266 226894
rect 333822 226338 333854 226894
rect 333234 190894 333854 226338
rect 333234 190338 333266 190894
rect 333822 190338 333854 190894
rect 333234 154894 333854 190338
rect 333234 154338 333266 154894
rect 333822 154338 333854 154894
rect 333234 118894 333854 154338
rect 333234 118338 333266 118894
rect 333822 118338 333854 118894
rect 333234 82894 333854 118338
rect 333234 82338 333266 82894
rect 333822 82338 333854 82894
rect 333234 46894 333854 82338
rect 333234 46338 333266 46894
rect 333822 46338 333854 46894
rect 333234 10894 333854 46338
rect 333234 10338 333266 10894
rect 333822 10338 333854 10894
rect 333234 -4186 333854 10338
rect 333234 -4742 333266 -4186
rect 333822 -4742 333854 -4186
rect 333234 -5734 333854 -4742
rect 336954 302614 337574 336000
rect 336954 302058 336986 302614
rect 337542 302058 337574 302614
rect 336954 266614 337574 302058
rect 336954 266058 336986 266614
rect 337542 266058 337574 266614
rect 336954 230614 337574 266058
rect 336954 230058 336986 230614
rect 337542 230058 337574 230614
rect 336954 194614 337574 230058
rect 336954 194058 336986 194614
rect 337542 194058 337574 194614
rect 336954 158614 337574 194058
rect 336954 158058 336986 158614
rect 337542 158058 337574 158614
rect 336954 122614 337574 158058
rect 336954 122058 336986 122614
rect 337542 122058 337574 122614
rect 336954 86614 337574 122058
rect 336954 86058 336986 86614
rect 337542 86058 337574 86614
rect 336954 50614 337574 86058
rect 336954 50058 336986 50614
rect 337542 50058 337574 50614
rect 336954 14614 337574 50058
rect 336954 14058 336986 14614
rect 337542 14058 337574 14614
rect 318954 -7622 318986 -7066
rect 319542 -7622 319574 -7066
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 309454 344414 338000
rect 343794 308898 343826 309454
rect 344382 308898 344414 309454
rect 343794 273454 344414 308898
rect 343794 272898 343826 273454
rect 344382 272898 344414 273454
rect 343794 237454 344414 272898
rect 343794 236898 343826 237454
rect 344382 236898 344414 237454
rect 343794 201454 344414 236898
rect 343794 200898 343826 201454
rect 344382 200898 344414 201454
rect 343794 165454 344414 200898
rect 343794 164898 343826 165454
rect 344382 164898 344414 165454
rect 343794 129454 344414 164898
rect 343794 128898 343826 129454
rect 344382 128898 344414 129454
rect 343794 93454 344414 128898
rect 343794 92898 343826 93454
rect 344382 92898 344414 93454
rect 343794 57454 344414 92898
rect 343794 56898 343826 57454
rect 344382 56898 344414 57454
rect 343794 21454 344414 56898
rect 343794 20898 343826 21454
rect 344382 20898 344414 21454
rect 343794 -1306 344414 20898
rect 343794 -1862 343826 -1306
rect 344382 -1862 344414 -1306
rect 343794 -1894 344414 -1862
rect 347514 313174 348134 336000
rect 347514 312618 347546 313174
rect 348102 312618 348134 313174
rect 347514 277174 348134 312618
rect 347514 276618 347546 277174
rect 348102 276618 348134 277174
rect 347514 241174 348134 276618
rect 347514 240618 347546 241174
rect 348102 240618 348134 241174
rect 347514 205174 348134 240618
rect 347514 204618 347546 205174
rect 348102 204618 348134 205174
rect 347514 169174 348134 204618
rect 347514 168618 347546 169174
rect 348102 168618 348134 169174
rect 347514 133174 348134 168618
rect 347514 132618 347546 133174
rect 348102 132618 348134 133174
rect 347514 97174 348134 132618
rect 347514 96618 347546 97174
rect 348102 96618 348134 97174
rect 347514 61174 348134 96618
rect 347514 60618 347546 61174
rect 348102 60618 348134 61174
rect 347514 25174 348134 60618
rect 347514 24618 347546 25174
rect 348102 24618 348134 25174
rect 347514 -3226 348134 24618
rect 347514 -3782 347546 -3226
rect 348102 -3782 348134 -3226
rect 347514 -3814 348134 -3782
rect 351234 316894 351854 336000
rect 351234 316338 351266 316894
rect 351822 316338 351854 316894
rect 351234 280894 351854 316338
rect 351234 280338 351266 280894
rect 351822 280338 351854 280894
rect 351234 244894 351854 280338
rect 351234 244338 351266 244894
rect 351822 244338 351854 244894
rect 351234 208894 351854 244338
rect 351234 208338 351266 208894
rect 351822 208338 351854 208894
rect 351234 172894 351854 208338
rect 351234 172338 351266 172894
rect 351822 172338 351854 172894
rect 351234 136894 351854 172338
rect 351234 136338 351266 136894
rect 351822 136338 351854 136894
rect 351234 100894 351854 136338
rect 351234 100338 351266 100894
rect 351822 100338 351854 100894
rect 351234 64894 351854 100338
rect 351234 64338 351266 64894
rect 351822 64338 351854 64894
rect 351234 28894 351854 64338
rect 351234 28338 351266 28894
rect 351822 28338 351854 28894
rect 351234 -5146 351854 28338
rect 351234 -5702 351266 -5146
rect 351822 -5702 351854 -5146
rect 351234 -5734 351854 -5702
rect 354954 320614 355574 336000
rect 354954 320058 354986 320614
rect 355542 320058 355574 320614
rect 354954 284614 355574 320058
rect 354954 284058 354986 284614
rect 355542 284058 355574 284614
rect 354954 248614 355574 284058
rect 354954 248058 354986 248614
rect 355542 248058 355574 248614
rect 354954 212614 355574 248058
rect 354954 212058 354986 212614
rect 355542 212058 355574 212614
rect 354954 176614 355574 212058
rect 354954 176058 354986 176614
rect 355542 176058 355574 176614
rect 354954 140614 355574 176058
rect 354954 140058 354986 140614
rect 355542 140058 355574 140614
rect 354954 104614 355574 140058
rect 354954 104058 354986 104614
rect 355542 104058 355574 104614
rect 354954 68614 355574 104058
rect 354954 68058 354986 68614
rect 355542 68058 355574 68614
rect 354954 32614 355574 68058
rect 354954 32058 354986 32614
rect 355542 32058 355574 32614
rect 336954 -6662 336986 -6106
rect 337542 -6662 337574 -6106
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 327454 362414 338000
rect 361794 326898 361826 327454
rect 362382 326898 362414 327454
rect 361794 291454 362414 326898
rect 361794 290898 361826 291454
rect 362382 290898 362414 291454
rect 361794 255454 362414 290898
rect 361794 254898 361826 255454
rect 362382 254898 362414 255454
rect 361794 219454 362414 254898
rect 361794 218898 361826 219454
rect 362382 218898 362414 219454
rect 361794 183454 362414 218898
rect 361794 182898 361826 183454
rect 362382 182898 362414 183454
rect 361794 147454 362414 182898
rect 361794 146898 361826 147454
rect 362382 146898 362414 147454
rect 361794 111454 362414 146898
rect 361794 110898 361826 111454
rect 362382 110898 362414 111454
rect 361794 75454 362414 110898
rect 361794 74898 361826 75454
rect 362382 74898 362414 75454
rect 361794 39454 362414 74898
rect 361794 38898 361826 39454
rect 362382 38898 362414 39454
rect 361794 3454 362414 38898
rect 361794 2898 361826 3454
rect 362382 2898 362414 3454
rect 361794 -346 362414 2898
rect 361794 -902 361826 -346
rect 362382 -902 362414 -346
rect 361794 -1894 362414 -902
rect 365514 331174 366134 336000
rect 365514 330618 365546 331174
rect 366102 330618 366134 331174
rect 365514 295174 366134 330618
rect 365514 294618 365546 295174
rect 366102 294618 366134 295174
rect 365514 259174 366134 294618
rect 365514 258618 365546 259174
rect 366102 258618 366134 259174
rect 365514 223174 366134 258618
rect 365514 222618 365546 223174
rect 366102 222618 366134 223174
rect 365514 187174 366134 222618
rect 365514 186618 365546 187174
rect 366102 186618 366134 187174
rect 365514 151174 366134 186618
rect 365514 150618 365546 151174
rect 366102 150618 366134 151174
rect 365514 115174 366134 150618
rect 365514 114618 365546 115174
rect 366102 114618 366134 115174
rect 365514 79174 366134 114618
rect 365514 78618 365546 79174
rect 366102 78618 366134 79174
rect 365514 43174 366134 78618
rect 365514 42618 365546 43174
rect 366102 42618 366134 43174
rect 365514 7174 366134 42618
rect 365514 6618 365546 7174
rect 366102 6618 366134 7174
rect 365514 -2266 366134 6618
rect 365514 -2822 365546 -2266
rect 366102 -2822 366134 -2266
rect 365514 -3814 366134 -2822
rect 369234 334894 369854 336000
rect 369234 334338 369266 334894
rect 369822 334338 369854 334894
rect 369234 298894 369854 334338
rect 369234 298338 369266 298894
rect 369822 298338 369854 298894
rect 369234 262894 369854 298338
rect 369234 262338 369266 262894
rect 369822 262338 369854 262894
rect 369234 226894 369854 262338
rect 369234 226338 369266 226894
rect 369822 226338 369854 226894
rect 369234 190894 369854 226338
rect 369234 190338 369266 190894
rect 369822 190338 369854 190894
rect 369234 154894 369854 190338
rect 369234 154338 369266 154894
rect 369822 154338 369854 154894
rect 369234 118894 369854 154338
rect 369234 118338 369266 118894
rect 369822 118338 369854 118894
rect 369234 82894 369854 118338
rect 369234 82338 369266 82894
rect 369822 82338 369854 82894
rect 369234 46894 369854 82338
rect 369234 46338 369266 46894
rect 369822 46338 369854 46894
rect 369234 10894 369854 46338
rect 369234 10338 369266 10894
rect 369822 10338 369854 10894
rect 369234 -4186 369854 10338
rect 369234 -4742 369266 -4186
rect 369822 -4742 369854 -4186
rect 369234 -5734 369854 -4742
rect 372954 302614 373574 336000
rect 372954 302058 372986 302614
rect 373542 302058 373574 302614
rect 372954 266614 373574 302058
rect 372954 266058 372986 266614
rect 373542 266058 373574 266614
rect 372954 230614 373574 266058
rect 372954 230058 372986 230614
rect 373542 230058 373574 230614
rect 372954 194614 373574 230058
rect 372954 194058 372986 194614
rect 373542 194058 373574 194614
rect 372954 158614 373574 194058
rect 372954 158058 372986 158614
rect 373542 158058 373574 158614
rect 372954 122614 373574 158058
rect 372954 122058 372986 122614
rect 373542 122058 373574 122614
rect 372954 86614 373574 122058
rect 372954 86058 372986 86614
rect 373542 86058 373574 86614
rect 372954 50614 373574 86058
rect 372954 50058 372986 50614
rect 373542 50058 373574 50614
rect 372954 14614 373574 50058
rect 372954 14058 372986 14614
rect 373542 14058 373574 14614
rect 354954 -7622 354986 -7066
rect 355542 -7622 355574 -7066
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 309454 380414 338000
rect 382230 320109 382290 457267
rect 382227 320108 382293 320109
rect 382227 320044 382228 320108
rect 382292 320044 382293 320108
rect 382227 320043 382293 320044
rect 379794 308898 379826 309454
rect 380382 308898 380414 309454
rect 379794 273454 380414 308898
rect 379794 272898 379826 273454
rect 380382 272898 380414 273454
rect 379794 237454 380414 272898
rect 379794 236898 379826 237454
rect 380382 236898 380414 237454
rect 379794 201454 380414 236898
rect 379794 200898 379826 201454
rect 380382 200898 380414 201454
rect 379794 165454 380414 200898
rect 379794 164898 379826 165454
rect 380382 164898 380414 165454
rect 379794 129454 380414 164898
rect 379794 128898 379826 129454
rect 380382 128898 380414 129454
rect 379794 93454 380414 128898
rect 379794 92898 379826 93454
rect 380382 92898 380414 93454
rect 379794 57454 380414 92898
rect 379794 56898 379826 57454
rect 380382 56898 380414 57454
rect 379794 21454 380414 56898
rect 379794 20898 379826 21454
rect 380382 20898 380414 21454
rect 379794 -1306 380414 20898
rect 379794 -1862 379826 -1306
rect 380382 -1862 380414 -1306
rect 379794 -1894 380414 -1862
rect 383514 313174 384134 336000
rect 383514 312618 383546 313174
rect 384102 312618 384134 313174
rect 383514 277174 384134 312618
rect 384254 293861 384314 457267
rect 384990 306373 385050 457267
rect 384987 306372 385053 306373
rect 384987 306308 384988 306372
rect 385052 306308 385053 306372
rect 384987 306307 385053 306308
rect 384251 293860 384317 293861
rect 384251 293796 384252 293860
rect 384316 293796 384317 293860
rect 384251 293795 384317 293796
rect 383514 276618 383546 277174
rect 384102 276618 384134 277174
rect 383514 241174 384134 276618
rect 386462 267749 386522 457267
rect 387234 316894 387854 336000
rect 387234 316338 387266 316894
rect 387822 316338 387854 316894
rect 387234 280894 387854 316338
rect 387234 280338 387266 280894
rect 387822 280338 387854 280894
rect 386459 267748 386525 267749
rect 386459 267684 386460 267748
rect 386524 267684 386525 267748
rect 386459 267683 386525 267684
rect 383514 240618 383546 241174
rect 384102 240618 384134 241174
rect 383514 205174 384134 240618
rect 383514 204618 383546 205174
rect 384102 204618 384134 205174
rect 383514 169174 384134 204618
rect 383514 168618 383546 169174
rect 384102 168618 384134 169174
rect 383514 133174 384134 168618
rect 383514 132618 383546 133174
rect 384102 132618 384134 133174
rect 383514 97174 384134 132618
rect 383514 96618 383546 97174
rect 384102 96618 384134 97174
rect 383514 61174 384134 96618
rect 383514 60618 383546 61174
rect 384102 60618 384134 61174
rect 383514 25174 384134 60618
rect 383514 24618 383546 25174
rect 384102 24618 384134 25174
rect 383514 -3226 384134 24618
rect 383514 -3782 383546 -3226
rect 384102 -3782 384134 -3226
rect 383514 -3814 384134 -3782
rect 387234 244894 387854 280338
rect 387934 248430 387994 457267
rect 389222 255237 389282 457267
rect 392808 435454 393128 435486
rect 392808 435218 392850 435454
rect 393086 435218 393128 435454
rect 392808 435134 393128 435218
rect 392808 434898 392850 435134
rect 393086 434898 393128 435134
rect 392808 434866 393128 434898
rect 392808 399454 393128 399486
rect 392808 399218 392850 399454
rect 393086 399218 393128 399454
rect 392808 399134 393128 399218
rect 392808 398898 392850 399134
rect 393086 398898 393128 399134
rect 392808 398866 393128 398898
rect 392808 363454 393128 363486
rect 392808 363218 392850 363454
rect 393086 363218 393128 363454
rect 392808 363134 393128 363218
rect 392808 362898 392850 363134
rect 393086 362898 393128 363134
rect 392808 362866 393128 362898
rect 393454 339690 393514 457267
rect 393086 339630 393514 339690
rect 390954 320614 391574 336000
rect 390954 320058 390986 320614
rect 391542 320058 391574 320614
rect 390954 284614 391574 320058
rect 390954 284058 390986 284614
rect 391542 284058 391574 284614
rect 389219 255236 389285 255237
rect 389219 255172 389220 255236
rect 389284 255172 389285 255236
rect 389219 255171 389285 255172
rect 390954 248614 391574 284058
rect 387934 248370 388178 248430
rect 387234 244338 387266 244894
rect 387822 244338 387854 244894
rect 387234 208894 387854 244338
rect 388118 241501 388178 248370
rect 390954 248058 390986 248614
rect 391542 248058 391574 248614
rect 388115 241500 388181 241501
rect 388115 241436 388116 241500
rect 388180 241436 388181 241500
rect 388115 241435 388181 241436
rect 387234 208338 387266 208894
rect 387822 208338 387854 208894
rect 387234 172894 387854 208338
rect 387234 172338 387266 172894
rect 387822 172338 387854 172894
rect 387234 136894 387854 172338
rect 387234 136338 387266 136894
rect 387822 136338 387854 136894
rect 387234 100894 387854 136338
rect 387234 100338 387266 100894
rect 387822 100338 387854 100894
rect 387234 64894 387854 100338
rect 387234 64338 387266 64894
rect 387822 64338 387854 64894
rect 387234 28894 387854 64338
rect 387234 28338 387266 28894
rect 387822 28338 387854 28894
rect 387234 -5146 387854 28338
rect 387234 -5702 387266 -5146
rect 387822 -5702 387854 -5146
rect 387234 -5734 387854 -5702
rect 390954 212614 391574 248058
rect 390954 212058 390986 212614
rect 391542 212058 391574 212614
rect 390954 176614 391574 212058
rect 393086 189005 393146 339630
rect 394742 202877 394802 457267
rect 394739 202876 394805 202877
rect 394739 202812 394740 202876
rect 394804 202812 394805 202876
rect 394739 202811 394805 202812
rect 393083 189004 393149 189005
rect 393083 188940 393084 189004
rect 393148 188940 393149 189004
rect 393083 188939 393149 188940
rect 390954 176058 390986 176614
rect 391542 176058 391574 176614
rect 390954 140614 391574 176058
rect 396214 164117 396274 457267
rect 396211 164116 396277 164117
rect 396211 164052 396212 164116
rect 396276 164052 396277 164116
rect 396211 164051 396277 164052
rect 390954 140058 390986 140614
rect 391542 140058 391574 140614
rect 390954 104614 391574 140058
rect 397502 138005 397562 457267
rect 397794 327454 398414 338000
rect 397794 326898 397826 327454
rect 398382 326898 398414 327454
rect 397794 291454 398414 326898
rect 397794 290898 397826 291454
rect 398382 290898 398414 291454
rect 397794 255454 398414 290898
rect 397794 254898 397826 255454
rect 398382 254898 398414 255454
rect 397794 219454 398414 254898
rect 397794 218898 397826 219454
rect 398382 218898 398414 219454
rect 397794 183454 398414 218898
rect 397794 182898 397826 183454
rect 398382 182898 398414 183454
rect 397794 147454 398414 182898
rect 398790 150381 398850 457267
rect 398787 150380 398853 150381
rect 398787 150316 398788 150380
rect 398852 150316 398853 150380
rect 398787 150315 398853 150316
rect 397794 146898 397826 147454
rect 398382 146898 398414 147454
rect 397499 138004 397565 138005
rect 397499 137940 397500 138004
rect 397564 137940 397565 138004
rect 397499 137939 397565 137940
rect 390954 104058 390986 104614
rect 391542 104058 391574 104614
rect 390954 68614 391574 104058
rect 390954 68058 390986 68614
rect 391542 68058 391574 68614
rect 390954 32614 391574 68058
rect 390954 32058 390986 32614
rect 391542 32058 391574 32614
rect 372954 -6662 372986 -6106
rect 373542 -6662 373574 -6106
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 111454 398414 146898
rect 400262 111757 400322 457267
rect 401514 331174 402134 336000
rect 401514 330618 401546 331174
rect 402102 330618 402134 331174
rect 401514 295174 402134 330618
rect 401514 294618 401546 295174
rect 402102 294618 402134 295174
rect 401514 259174 402134 294618
rect 401514 258618 401546 259174
rect 402102 258618 402134 259174
rect 401514 223174 402134 258618
rect 401514 222618 401546 223174
rect 402102 222618 402134 223174
rect 401514 187174 402134 222618
rect 401514 186618 401546 187174
rect 402102 186618 402134 187174
rect 401514 151174 402134 186618
rect 401514 150618 401546 151174
rect 402102 150618 402134 151174
rect 401514 115174 402134 150618
rect 401514 114618 401546 115174
rect 402102 114618 402134 115174
rect 400259 111756 400325 111757
rect 400259 111692 400260 111756
rect 400324 111692 400325 111756
rect 400259 111691 400325 111692
rect 397794 110898 397826 111454
rect 398382 110898 398414 111454
rect 397794 75454 398414 110898
rect 397794 74898 397826 75454
rect 398382 74898 398414 75454
rect 397794 39454 398414 74898
rect 397794 38898 397826 39454
rect 398382 38898 398414 39454
rect 397794 3454 398414 38898
rect 397794 2898 397826 3454
rect 398382 2898 398414 3454
rect 397794 -346 398414 2898
rect 397794 -902 397826 -346
rect 398382 -902 398414 -346
rect 397794 -1894 398414 -902
rect 401514 79174 402134 114618
rect 403022 85509 403082 457267
rect 404310 97885 404370 457267
rect 405234 334894 405854 336000
rect 405234 334338 405266 334894
rect 405822 334338 405854 334894
rect 405234 298894 405854 334338
rect 405234 298338 405266 298894
rect 405822 298338 405854 298894
rect 405234 262894 405854 298338
rect 405234 262338 405266 262894
rect 405822 262338 405854 262894
rect 405234 226894 405854 262338
rect 405234 226338 405266 226894
rect 405822 226338 405854 226894
rect 405234 190894 405854 226338
rect 405234 190338 405266 190894
rect 405822 190338 405854 190894
rect 405234 154894 405854 190338
rect 405234 154338 405266 154894
rect 405822 154338 405854 154894
rect 405234 118894 405854 154338
rect 405234 118338 405266 118894
rect 405822 118338 405854 118894
rect 404307 97884 404373 97885
rect 404307 97820 404308 97884
rect 404372 97820 404373 97884
rect 404307 97819 404373 97820
rect 403019 85508 403085 85509
rect 403019 85444 403020 85508
rect 403084 85444 403085 85508
rect 403019 85443 403085 85444
rect 401514 78618 401546 79174
rect 402102 78618 402134 79174
rect 401514 43174 402134 78618
rect 401514 42618 401546 43174
rect 402102 42618 402134 43174
rect 401514 7174 402134 42618
rect 401514 6618 401546 7174
rect 402102 6618 402134 7174
rect 401514 -2266 402134 6618
rect 401514 -2822 401546 -2266
rect 402102 -2822 402134 -2266
rect 401514 -3814 402134 -2822
rect 405234 82894 405854 118338
rect 405234 82338 405266 82894
rect 405822 82338 405854 82894
rect 405234 46894 405854 82338
rect 405966 71773 406026 457267
rect 408168 453454 408488 453486
rect 408168 453218 408210 453454
rect 408446 453218 408488 453454
rect 408168 453134 408488 453218
rect 408168 452898 408210 453134
rect 408446 452898 408488 453134
rect 408168 452866 408488 452898
rect 408168 417454 408488 417486
rect 408168 417218 408210 417454
rect 408446 417218 408488 417454
rect 408168 417134 408488 417218
rect 408168 416898 408210 417134
rect 408446 416898 408488 417134
rect 408168 416866 408488 416898
rect 408168 381454 408488 381486
rect 408168 381218 408210 381454
rect 408446 381218 408488 381454
rect 408168 381134 408488 381218
rect 408168 380898 408210 381134
rect 408446 380898 408488 381134
rect 408168 380866 408488 380898
rect 408168 345454 408488 345486
rect 408168 345218 408210 345454
rect 408446 345218 408488 345454
rect 408168 345134 408488 345218
rect 408168 344898 408210 345134
rect 408446 344898 408488 345134
rect 408168 344866 408488 344898
rect 405963 71772 406029 71773
rect 405963 71708 405964 71772
rect 406028 71708 406029 71772
rect 405963 71707 406029 71708
rect 408726 59261 408786 457267
rect 408954 302614 409574 336000
rect 408954 302058 408986 302614
rect 409542 302058 409574 302614
rect 408954 266614 409574 302058
rect 408954 266058 408986 266614
rect 409542 266058 409574 266614
rect 408954 230614 409574 266058
rect 408954 230058 408986 230614
rect 409542 230058 409574 230614
rect 408954 194614 409574 230058
rect 408954 194058 408986 194614
rect 409542 194058 409574 194614
rect 408954 158614 409574 194058
rect 408954 158058 408986 158614
rect 409542 158058 409574 158614
rect 408954 122614 409574 158058
rect 408954 122058 408986 122614
rect 409542 122058 409574 122614
rect 408954 86614 409574 122058
rect 408954 86058 408986 86614
rect 409542 86058 409574 86614
rect 408723 59260 408789 59261
rect 408723 59196 408724 59260
rect 408788 59196 408789 59260
rect 408723 59195 408789 59196
rect 405234 46338 405266 46894
rect 405822 46338 405854 46894
rect 405234 10894 405854 46338
rect 405234 10338 405266 10894
rect 405822 10338 405854 10894
rect 405234 -4186 405854 10338
rect 405234 -4742 405266 -4186
rect 405822 -4742 405854 -4186
rect 405234 -5734 405854 -4742
rect 408954 50614 409574 86058
rect 408954 50058 408986 50614
rect 409542 50058 409574 50614
rect 408954 14614 409574 50058
rect 409830 33149 409890 457267
rect 409827 33148 409893 33149
rect 409827 33084 409828 33148
rect 409892 33084 409893 33148
rect 409827 33083 409893 33084
rect 408954 14058 408986 14614
rect 409542 14058 409574 14614
rect 390954 -7622 390986 -7066
rect 391542 -7622 391574 -7066
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 411302 6901 411362 457267
rect 415794 453454 416414 488898
rect 415794 452898 415826 453454
rect 416382 452898 416414 453454
rect 415794 417454 416414 452898
rect 415794 416898 415826 417454
rect 416382 416898 416414 417454
rect 415794 381454 416414 416898
rect 415794 380898 415826 381454
rect 416382 380898 416414 381454
rect 415794 345454 416414 380898
rect 415794 344898 415826 345454
rect 416382 344898 416414 345454
rect 415794 309454 416414 344898
rect 415794 308898 415826 309454
rect 416382 308898 416414 309454
rect 415794 273454 416414 308898
rect 415794 272898 415826 273454
rect 416382 272898 416414 273454
rect 415794 237454 416414 272898
rect 415794 236898 415826 237454
rect 416382 236898 416414 237454
rect 415794 201454 416414 236898
rect 415794 200898 415826 201454
rect 416382 200898 416414 201454
rect 415794 165454 416414 200898
rect 415794 164898 415826 165454
rect 416382 164898 416414 165454
rect 415794 129454 416414 164898
rect 415794 128898 415826 129454
rect 416382 128898 416414 129454
rect 415794 93454 416414 128898
rect 415794 92898 415826 93454
rect 416382 92898 416414 93454
rect 415794 57454 416414 92898
rect 415794 56898 415826 57454
rect 416382 56898 416414 57454
rect 415794 21454 416414 56898
rect 415794 20898 415826 21454
rect 416382 20898 416414 21454
rect 411299 6900 411365 6901
rect 411299 6836 411300 6900
rect 411364 6836 411365 6900
rect 411299 6835 411365 6836
rect 415794 -1306 416414 20898
rect 415794 -1862 415826 -1306
rect 416382 -1862 416414 -1306
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672618 419546 673174
rect 420102 672618 420134 673174
rect 419514 637174 420134 672618
rect 419514 636618 419546 637174
rect 420102 636618 420134 637174
rect 419514 601174 420134 636618
rect 419514 600618 419546 601174
rect 420102 600618 420134 601174
rect 419514 565174 420134 600618
rect 419514 564618 419546 565174
rect 420102 564618 420134 565174
rect 419514 529174 420134 564618
rect 419514 528618 419546 529174
rect 420102 528618 420134 529174
rect 419514 493174 420134 528618
rect 419514 492618 419546 493174
rect 420102 492618 420134 493174
rect 419514 457174 420134 492618
rect 419514 456618 419546 457174
rect 420102 456618 420134 457174
rect 419514 421174 420134 456618
rect 419514 420618 419546 421174
rect 420102 420618 420134 421174
rect 419514 385174 420134 420618
rect 419514 384618 419546 385174
rect 420102 384618 420134 385174
rect 419514 349174 420134 384618
rect 419514 348618 419546 349174
rect 420102 348618 420134 349174
rect 419514 313174 420134 348618
rect 419514 312618 419546 313174
rect 420102 312618 420134 313174
rect 419514 277174 420134 312618
rect 419514 276618 419546 277174
rect 420102 276618 420134 277174
rect 419514 241174 420134 276618
rect 419514 240618 419546 241174
rect 420102 240618 420134 241174
rect 419514 205174 420134 240618
rect 419514 204618 419546 205174
rect 420102 204618 420134 205174
rect 419514 169174 420134 204618
rect 419514 168618 419546 169174
rect 420102 168618 420134 169174
rect 419514 133174 420134 168618
rect 419514 132618 419546 133174
rect 420102 132618 420134 133174
rect 419514 97174 420134 132618
rect 419514 96618 419546 97174
rect 420102 96618 420134 97174
rect 419514 61174 420134 96618
rect 419514 60618 419546 61174
rect 420102 60618 420134 61174
rect 419514 25174 420134 60618
rect 419514 24618 419546 25174
rect 420102 24618 420134 25174
rect 419514 -3226 420134 24618
rect 419514 -3782 419546 -3226
rect 420102 -3782 420134 -3226
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676338 423266 676894
rect 423822 676338 423854 676894
rect 423234 640894 423854 676338
rect 423234 640338 423266 640894
rect 423822 640338 423854 640894
rect 423234 604894 423854 640338
rect 423234 604338 423266 604894
rect 423822 604338 423854 604894
rect 423234 568894 423854 604338
rect 423234 568338 423266 568894
rect 423822 568338 423854 568894
rect 423234 532894 423854 568338
rect 423234 532338 423266 532894
rect 423822 532338 423854 532894
rect 423234 496894 423854 532338
rect 423234 496338 423266 496894
rect 423822 496338 423854 496894
rect 423234 460894 423854 496338
rect 423234 460338 423266 460894
rect 423822 460338 423854 460894
rect 423234 424894 423854 460338
rect 423234 424338 423266 424894
rect 423822 424338 423854 424894
rect 423234 388894 423854 424338
rect 423234 388338 423266 388894
rect 423822 388338 423854 388894
rect 423234 352894 423854 388338
rect 423234 352338 423266 352894
rect 423822 352338 423854 352894
rect 423234 316894 423854 352338
rect 423234 316338 423266 316894
rect 423822 316338 423854 316894
rect 423234 280894 423854 316338
rect 423234 280338 423266 280894
rect 423822 280338 423854 280894
rect 423234 244894 423854 280338
rect 423234 244338 423266 244894
rect 423822 244338 423854 244894
rect 423234 208894 423854 244338
rect 423234 208338 423266 208894
rect 423822 208338 423854 208894
rect 423234 172894 423854 208338
rect 423234 172338 423266 172894
rect 423822 172338 423854 172894
rect 423234 136894 423854 172338
rect 423234 136338 423266 136894
rect 423822 136338 423854 136894
rect 423234 100894 423854 136338
rect 423234 100338 423266 100894
rect 423822 100338 423854 100894
rect 423234 64894 423854 100338
rect 423234 64338 423266 64894
rect 423822 64338 423854 64894
rect 423234 28894 423854 64338
rect 423234 28338 423266 28894
rect 423822 28338 423854 28894
rect 423234 -5146 423854 28338
rect 423234 -5702 423266 -5146
rect 423822 -5702 423854 -5146
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710042 444986 710598
rect 445542 710042 445574 710598
rect 441234 708678 441854 709670
rect 441234 708122 441266 708678
rect 441822 708122 441854 708678
rect 437514 706758 438134 707750
rect 437514 706202 437546 706758
rect 438102 706202 438134 706758
rect 426954 680058 426986 680614
rect 427542 680058 427574 680614
rect 426954 644614 427574 680058
rect 426954 644058 426986 644614
rect 427542 644058 427574 644614
rect 426954 608614 427574 644058
rect 426954 608058 426986 608614
rect 427542 608058 427574 608614
rect 426954 572614 427574 608058
rect 426954 572058 426986 572614
rect 427542 572058 427574 572614
rect 426954 536614 427574 572058
rect 426954 536058 426986 536614
rect 427542 536058 427574 536614
rect 426954 500614 427574 536058
rect 426954 500058 426986 500614
rect 427542 500058 427574 500614
rect 426954 464614 427574 500058
rect 426954 464058 426986 464614
rect 427542 464058 427574 464614
rect 426954 428614 427574 464058
rect 426954 428058 426986 428614
rect 427542 428058 427574 428614
rect 426954 392614 427574 428058
rect 426954 392058 426986 392614
rect 427542 392058 427574 392614
rect 426954 356614 427574 392058
rect 426954 356058 426986 356614
rect 427542 356058 427574 356614
rect 426954 320614 427574 356058
rect 426954 320058 426986 320614
rect 427542 320058 427574 320614
rect 426954 284614 427574 320058
rect 426954 284058 426986 284614
rect 427542 284058 427574 284614
rect 426954 248614 427574 284058
rect 426954 248058 426986 248614
rect 427542 248058 427574 248614
rect 426954 212614 427574 248058
rect 426954 212058 426986 212614
rect 427542 212058 427574 212614
rect 426954 176614 427574 212058
rect 426954 176058 426986 176614
rect 427542 176058 427574 176614
rect 426954 140614 427574 176058
rect 426954 140058 426986 140614
rect 427542 140058 427574 140614
rect 426954 104614 427574 140058
rect 426954 104058 426986 104614
rect 427542 104058 427574 104614
rect 426954 68614 427574 104058
rect 426954 68058 426986 68614
rect 427542 68058 427574 68614
rect 426954 32614 427574 68058
rect 426954 32058 426986 32614
rect 427542 32058 427574 32614
rect 408954 -6662 408986 -6106
rect 409542 -6662 409574 -6106
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704282 433826 704838
rect 434382 704282 434414 704838
rect 433794 687454 434414 704282
rect 433794 686898 433826 687454
rect 434382 686898 434414 687454
rect 433794 651454 434414 686898
rect 433794 650898 433826 651454
rect 434382 650898 434414 651454
rect 433794 615454 434414 650898
rect 433794 614898 433826 615454
rect 434382 614898 434414 615454
rect 433794 579454 434414 614898
rect 433794 578898 433826 579454
rect 434382 578898 434414 579454
rect 433794 543454 434414 578898
rect 433794 542898 433826 543454
rect 434382 542898 434414 543454
rect 433794 507454 434414 542898
rect 433794 506898 433826 507454
rect 434382 506898 434414 507454
rect 433794 471454 434414 506898
rect 433794 470898 433826 471454
rect 434382 470898 434414 471454
rect 433794 435454 434414 470898
rect 433794 434898 433826 435454
rect 434382 434898 434414 435454
rect 433794 399454 434414 434898
rect 433794 398898 433826 399454
rect 434382 398898 434414 399454
rect 433794 363454 434414 398898
rect 433794 362898 433826 363454
rect 434382 362898 434414 363454
rect 433794 327454 434414 362898
rect 433794 326898 433826 327454
rect 434382 326898 434414 327454
rect 433794 291454 434414 326898
rect 433794 290898 433826 291454
rect 434382 290898 434414 291454
rect 433794 255454 434414 290898
rect 433794 254898 433826 255454
rect 434382 254898 434414 255454
rect 433794 219454 434414 254898
rect 433794 218898 433826 219454
rect 434382 218898 434414 219454
rect 433794 183454 434414 218898
rect 433794 182898 433826 183454
rect 434382 182898 434414 183454
rect 433794 147454 434414 182898
rect 433794 146898 433826 147454
rect 434382 146898 434414 147454
rect 433794 111454 434414 146898
rect 433794 110898 433826 111454
rect 434382 110898 434414 111454
rect 433794 75454 434414 110898
rect 433794 74898 433826 75454
rect 434382 74898 434414 75454
rect 433794 39454 434414 74898
rect 433794 38898 433826 39454
rect 434382 38898 434414 39454
rect 433794 3454 434414 38898
rect 433794 2898 433826 3454
rect 434382 2898 434414 3454
rect 433794 -346 434414 2898
rect 433794 -902 433826 -346
rect 434382 -902 434414 -346
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690618 437546 691174
rect 438102 690618 438134 691174
rect 437514 655174 438134 690618
rect 437514 654618 437546 655174
rect 438102 654618 438134 655174
rect 437514 619174 438134 654618
rect 437514 618618 437546 619174
rect 438102 618618 438134 619174
rect 437514 583174 438134 618618
rect 437514 582618 437546 583174
rect 438102 582618 438134 583174
rect 437514 547174 438134 582618
rect 437514 546618 437546 547174
rect 438102 546618 438134 547174
rect 437514 511174 438134 546618
rect 437514 510618 437546 511174
rect 438102 510618 438134 511174
rect 437514 475174 438134 510618
rect 437514 474618 437546 475174
rect 438102 474618 438134 475174
rect 437514 439174 438134 474618
rect 437514 438618 437546 439174
rect 438102 438618 438134 439174
rect 437514 403174 438134 438618
rect 437514 402618 437546 403174
rect 438102 402618 438134 403174
rect 437514 367174 438134 402618
rect 437514 366618 437546 367174
rect 438102 366618 438134 367174
rect 437514 331174 438134 366618
rect 437514 330618 437546 331174
rect 438102 330618 438134 331174
rect 437514 295174 438134 330618
rect 437514 294618 437546 295174
rect 438102 294618 438134 295174
rect 437514 259174 438134 294618
rect 437514 258618 437546 259174
rect 438102 258618 438134 259174
rect 437514 223174 438134 258618
rect 437514 222618 437546 223174
rect 438102 222618 438134 223174
rect 437514 187174 438134 222618
rect 437514 186618 437546 187174
rect 438102 186618 438134 187174
rect 437514 151174 438134 186618
rect 437514 150618 437546 151174
rect 438102 150618 438134 151174
rect 437514 115174 438134 150618
rect 437514 114618 437546 115174
rect 438102 114618 438134 115174
rect 437514 79174 438134 114618
rect 437514 78618 437546 79174
rect 438102 78618 438134 79174
rect 437514 43174 438134 78618
rect 437514 42618 437546 43174
rect 438102 42618 438134 43174
rect 437514 7174 438134 42618
rect 437514 6618 437546 7174
rect 438102 6618 438134 7174
rect 437514 -2266 438134 6618
rect 437514 -2822 437546 -2266
rect 438102 -2822 438134 -2266
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694338 441266 694894
rect 441822 694338 441854 694894
rect 441234 658894 441854 694338
rect 441234 658338 441266 658894
rect 441822 658338 441854 658894
rect 441234 622894 441854 658338
rect 441234 622338 441266 622894
rect 441822 622338 441854 622894
rect 441234 586894 441854 622338
rect 441234 586338 441266 586894
rect 441822 586338 441854 586894
rect 441234 550894 441854 586338
rect 441234 550338 441266 550894
rect 441822 550338 441854 550894
rect 441234 514894 441854 550338
rect 441234 514338 441266 514894
rect 441822 514338 441854 514894
rect 441234 478894 441854 514338
rect 441234 478338 441266 478894
rect 441822 478338 441854 478894
rect 441234 442894 441854 478338
rect 441234 442338 441266 442894
rect 441822 442338 441854 442894
rect 441234 406894 441854 442338
rect 441234 406338 441266 406894
rect 441822 406338 441854 406894
rect 441234 370894 441854 406338
rect 441234 370338 441266 370894
rect 441822 370338 441854 370894
rect 441234 334894 441854 370338
rect 441234 334338 441266 334894
rect 441822 334338 441854 334894
rect 441234 298894 441854 334338
rect 441234 298338 441266 298894
rect 441822 298338 441854 298894
rect 441234 262894 441854 298338
rect 441234 262338 441266 262894
rect 441822 262338 441854 262894
rect 441234 226894 441854 262338
rect 441234 226338 441266 226894
rect 441822 226338 441854 226894
rect 441234 190894 441854 226338
rect 441234 190338 441266 190894
rect 441822 190338 441854 190894
rect 441234 154894 441854 190338
rect 441234 154338 441266 154894
rect 441822 154338 441854 154894
rect 441234 118894 441854 154338
rect 441234 118338 441266 118894
rect 441822 118338 441854 118894
rect 441234 82894 441854 118338
rect 441234 82338 441266 82894
rect 441822 82338 441854 82894
rect 441234 46894 441854 82338
rect 441234 46338 441266 46894
rect 441822 46338 441854 46894
rect 441234 10894 441854 46338
rect 441234 10338 441266 10894
rect 441822 10338 441854 10894
rect 441234 -4186 441854 10338
rect 441234 -4742 441266 -4186
rect 441822 -4742 441854 -4186
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711002 462986 711558
rect 463542 711002 463574 711558
rect 459234 709638 459854 709670
rect 459234 709082 459266 709638
rect 459822 709082 459854 709638
rect 455514 707718 456134 707750
rect 455514 707162 455546 707718
rect 456102 707162 456134 707718
rect 444954 698058 444986 698614
rect 445542 698058 445574 698614
rect 444954 662614 445574 698058
rect 444954 662058 444986 662614
rect 445542 662058 445574 662614
rect 444954 626614 445574 662058
rect 444954 626058 444986 626614
rect 445542 626058 445574 626614
rect 444954 590614 445574 626058
rect 444954 590058 444986 590614
rect 445542 590058 445574 590614
rect 444954 554614 445574 590058
rect 444954 554058 444986 554614
rect 445542 554058 445574 554614
rect 444954 518614 445574 554058
rect 444954 518058 444986 518614
rect 445542 518058 445574 518614
rect 444954 482614 445574 518058
rect 444954 482058 444986 482614
rect 445542 482058 445574 482614
rect 444954 446614 445574 482058
rect 444954 446058 444986 446614
rect 445542 446058 445574 446614
rect 444954 410614 445574 446058
rect 444954 410058 444986 410614
rect 445542 410058 445574 410614
rect 444954 374614 445574 410058
rect 444954 374058 444986 374614
rect 445542 374058 445574 374614
rect 444954 338614 445574 374058
rect 444954 338058 444986 338614
rect 445542 338058 445574 338614
rect 444954 302614 445574 338058
rect 444954 302058 444986 302614
rect 445542 302058 445574 302614
rect 444954 266614 445574 302058
rect 444954 266058 444986 266614
rect 445542 266058 445574 266614
rect 444954 230614 445574 266058
rect 444954 230058 444986 230614
rect 445542 230058 445574 230614
rect 444954 194614 445574 230058
rect 444954 194058 444986 194614
rect 445542 194058 445574 194614
rect 444954 158614 445574 194058
rect 444954 158058 444986 158614
rect 445542 158058 445574 158614
rect 444954 122614 445574 158058
rect 444954 122058 444986 122614
rect 445542 122058 445574 122614
rect 444954 86614 445574 122058
rect 444954 86058 444986 86614
rect 445542 86058 445574 86614
rect 444954 50614 445574 86058
rect 444954 50058 444986 50614
rect 445542 50058 445574 50614
rect 444954 14614 445574 50058
rect 444954 14058 444986 14614
rect 445542 14058 445574 14614
rect 426954 -7622 426986 -7066
rect 427542 -7622 427574 -7066
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705242 451826 705798
rect 452382 705242 452414 705798
rect 451794 669454 452414 705242
rect 451794 668898 451826 669454
rect 452382 668898 452414 669454
rect 451794 633454 452414 668898
rect 451794 632898 451826 633454
rect 452382 632898 452414 633454
rect 451794 597454 452414 632898
rect 451794 596898 451826 597454
rect 452382 596898 452414 597454
rect 451794 561454 452414 596898
rect 451794 560898 451826 561454
rect 452382 560898 452414 561454
rect 451794 525454 452414 560898
rect 451794 524898 451826 525454
rect 452382 524898 452414 525454
rect 451794 489454 452414 524898
rect 451794 488898 451826 489454
rect 452382 488898 452414 489454
rect 451794 453454 452414 488898
rect 451794 452898 451826 453454
rect 452382 452898 452414 453454
rect 451794 417454 452414 452898
rect 451794 416898 451826 417454
rect 452382 416898 452414 417454
rect 451794 381454 452414 416898
rect 451794 380898 451826 381454
rect 452382 380898 452414 381454
rect 451794 345454 452414 380898
rect 451794 344898 451826 345454
rect 452382 344898 452414 345454
rect 451794 309454 452414 344898
rect 451794 308898 451826 309454
rect 452382 308898 452414 309454
rect 451794 273454 452414 308898
rect 451794 272898 451826 273454
rect 452382 272898 452414 273454
rect 451794 237454 452414 272898
rect 451794 236898 451826 237454
rect 452382 236898 452414 237454
rect 451794 201454 452414 236898
rect 451794 200898 451826 201454
rect 452382 200898 452414 201454
rect 451794 165454 452414 200898
rect 451794 164898 451826 165454
rect 452382 164898 452414 165454
rect 451794 129454 452414 164898
rect 451794 128898 451826 129454
rect 452382 128898 452414 129454
rect 451794 93454 452414 128898
rect 451794 92898 451826 93454
rect 452382 92898 452414 93454
rect 451794 57454 452414 92898
rect 451794 56898 451826 57454
rect 452382 56898 452414 57454
rect 451794 21454 452414 56898
rect 451794 20898 451826 21454
rect 452382 20898 452414 21454
rect 451794 -1306 452414 20898
rect 451794 -1862 451826 -1306
rect 452382 -1862 452414 -1306
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672618 455546 673174
rect 456102 672618 456134 673174
rect 455514 637174 456134 672618
rect 455514 636618 455546 637174
rect 456102 636618 456134 637174
rect 455514 601174 456134 636618
rect 455514 600618 455546 601174
rect 456102 600618 456134 601174
rect 455514 565174 456134 600618
rect 455514 564618 455546 565174
rect 456102 564618 456134 565174
rect 455514 529174 456134 564618
rect 455514 528618 455546 529174
rect 456102 528618 456134 529174
rect 455514 493174 456134 528618
rect 455514 492618 455546 493174
rect 456102 492618 456134 493174
rect 455514 457174 456134 492618
rect 455514 456618 455546 457174
rect 456102 456618 456134 457174
rect 455514 421174 456134 456618
rect 455514 420618 455546 421174
rect 456102 420618 456134 421174
rect 455514 385174 456134 420618
rect 455514 384618 455546 385174
rect 456102 384618 456134 385174
rect 455514 349174 456134 384618
rect 455514 348618 455546 349174
rect 456102 348618 456134 349174
rect 455514 313174 456134 348618
rect 455514 312618 455546 313174
rect 456102 312618 456134 313174
rect 455514 277174 456134 312618
rect 455514 276618 455546 277174
rect 456102 276618 456134 277174
rect 455514 241174 456134 276618
rect 455514 240618 455546 241174
rect 456102 240618 456134 241174
rect 455514 205174 456134 240618
rect 455514 204618 455546 205174
rect 456102 204618 456134 205174
rect 455514 169174 456134 204618
rect 455514 168618 455546 169174
rect 456102 168618 456134 169174
rect 455514 133174 456134 168618
rect 455514 132618 455546 133174
rect 456102 132618 456134 133174
rect 455514 97174 456134 132618
rect 455514 96618 455546 97174
rect 456102 96618 456134 97174
rect 455514 61174 456134 96618
rect 455514 60618 455546 61174
rect 456102 60618 456134 61174
rect 455514 25174 456134 60618
rect 455514 24618 455546 25174
rect 456102 24618 456134 25174
rect 455514 -3226 456134 24618
rect 455514 -3782 455546 -3226
rect 456102 -3782 456134 -3226
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676338 459266 676894
rect 459822 676338 459854 676894
rect 459234 640894 459854 676338
rect 459234 640338 459266 640894
rect 459822 640338 459854 640894
rect 459234 604894 459854 640338
rect 459234 604338 459266 604894
rect 459822 604338 459854 604894
rect 459234 568894 459854 604338
rect 459234 568338 459266 568894
rect 459822 568338 459854 568894
rect 459234 532894 459854 568338
rect 459234 532338 459266 532894
rect 459822 532338 459854 532894
rect 459234 496894 459854 532338
rect 459234 496338 459266 496894
rect 459822 496338 459854 496894
rect 459234 460894 459854 496338
rect 459234 460338 459266 460894
rect 459822 460338 459854 460894
rect 459234 424894 459854 460338
rect 459234 424338 459266 424894
rect 459822 424338 459854 424894
rect 459234 388894 459854 424338
rect 459234 388338 459266 388894
rect 459822 388338 459854 388894
rect 459234 352894 459854 388338
rect 459234 352338 459266 352894
rect 459822 352338 459854 352894
rect 459234 316894 459854 352338
rect 459234 316338 459266 316894
rect 459822 316338 459854 316894
rect 459234 280894 459854 316338
rect 459234 280338 459266 280894
rect 459822 280338 459854 280894
rect 459234 244894 459854 280338
rect 459234 244338 459266 244894
rect 459822 244338 459854 244894
rect 459234 208894 459854 244338
rect 459234 208338 459266 208894
rect 459822 208338 459854 208894
rect 459234 172894 459854 208338
rect 459234 172338 459266 172894
rect 459822 172338 459854 172894
rect 459234 136894 459854 172338
rect 459234 136338 459266 136894
rect 459822 136338 459854 136894
rect 459234 100894 459854 136338
rect 459234 100338 459266 100894
rect 459822 100338 459854 100894
rect 459234 64894 459854 100338
rect 459234 64338 459266 64894
rect 459822 64338 459854 64894
rect 459234 28894 459854 64338
rect 459234 28338 459266 28894
rect 459822 28338 459854 28894
rect 459234 -5146 459854 28338
rect 459234 -5702 459266 -5146
rect 459822 -5702 459854 -5146
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710042 480986 710598
rect 481542 710042 481574 710598
rect 477234 708678 477854 709670
rect 477234 708122 477266 708678
rect 477822 708122 477854 708678
rect 473514 706758 474134 707750
rect 473514 706202 473546 706758
rect 474102 706202 474134 706758
rect 462954 680058 462986 680614
rect 463542 680058 463574 680614
rect 462954 644614 463574 680058
rect 462954 644058 462986 644614
rect 463542 644058 463574 644614
rect 462954 608614 463574 644058
rect 462954 608058 462986 608614
rect 463542 608058 463574 608614
rect 462954 572614 463574 608058
rect 462954 572058 462986 572614
rect 463542 572058 463574 572614
rect 462954 536614 463574 572058
rect 462954 536058 462986 536614
rect 463542 536058 463574 536614
rect 462954 500614 463574 536058
rect 462954 500058 462986 500614
rect 463542 500058 463574 500614
rect 462954 464614 463574 500058
rect 462954 464058 462986 464614
rect 463542 464058 463574 464614
rect 462954 428614 463574 464058
rect 462954 428058 462986 428614
rect 463542 428058 463574 428614
rect 462954 392614 463574 428058
rect 462954 392058 462986 392614
rect 463542 392058 463574 392614
rect 462954 356614 463574 392058
rect 462954 356058 462986 356614
rect 463542 356058 463574 356614
rect 462954 320614 463574 356058
rect 462954 320058 462986 320614
rect 463542 320058 463574 320614
rect 462954 284614 463574 320058
rect 462954 284058 462986 284614
rect 463542 284058 463574 284614
rect 462954 248614 463574 284058
rect 462954 248058 462986 248614
rect 463542 248058 463574 248614
rect 462954 212614 463574 248058
rect 462954 212058 462986 212614
rect 463542 212058 463574 212614
rect 462954 176614 463574 212058
rect 462954 176058 462986 176614
rect 463542 176058 463574 176614
rect 462954 140614 463574 176058
rect 462954 140058 462986 140614
rect 463542 140058 463574 140614
rect 462954 104614 463574 140058
rect 462954 104058 462986 104614
rect 463542 104058 463574 104614
rect 462954 68614 463574 104058
rect 462954 68058 462986 68614
rect 463542 68058 463574 68614
rect 462954 32614 463574 68058
rect 462954 32058 462986 32614
rect 463542 32058 463574 32614
rect 444954 -6662 444986 -6106
rect 445542 -6662 445574 -6106
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704282 469826 704838
rect 470382 704282 470414 704838
rect 469794 687454 470414 704282
rect 469794 686898 469826 687454
rect 470382 686898 470414 687454
rect 469794 651454 470414 686898
rect 469794 650898 469826 651454
rect 470382 650898 470414 651454
rect 469794 615454 470414 650898
rect 469794 614898 469826 615454
rect 470382 614898 470414 615454
rect 469794 579454 470414 614898
rect 469794 578898 469826 579454
rect 470382 578898 470414 579454
rect 469794 543454 470414 578898
rect 469794 542898 469826 543454
rect 470382 542898 470414 543454
rect 469794 507454 470414 542898
rect 469794 506898 469826 507454
rect 470382 506898 470414 507454
rect 469794 471454 470414 506898
rect 469794 470898 469826 471454
rect 470382 470898 470414 471454
rect 469794 435454 470414 470898
rect 469794 434898 469826 435454
rect 470382 434898 470414 435454
rect 469794 399454 470414 434898
rect 469794 398898 469826 399454
rect 470382 398898 470414 399454
rect 469794 363454 470414 398898
rect 469794 362898 469826 363454
rect 470382 362898 470414 363454
rect 469794 327454 470414 362898
rect 469794 326898 469826 327454
rect 470382 326898 470414 327454
rect 469794 291454 470414 326898
rect 469794 290898 469826 291454
rect 470382 290898 470414 291454
rect 469794 255454 470414 290898
rect 469794 254898 469826 255454
rect 470382 254898 470414 255454
rect 469794 219454 470414 254898
rect 469794 218898 469826 219454
rect 470382 218898 470414 219454
rect 469794 183454 470414 218898
rect 469794 182898 469826 183454
rect 470382 182898 470414 183454
rect 469794 147454 470414 182898
rect 469794 146898 469826 147454
rect 470382 146898 470414 147454
rect 469794 111454 470414 146898
rect 469794 110898 469826 111454
rect 470382 110898 470414 111454
rect 469794 75454 470414 110898
rect 469794 74898 469826 75454
rect 470382 74898 470414 75454
rect 469794 39454 470414 74898
rect 469794 38898 469826 39454
rect 470382 38898 470414 39454
rect 469794 3454 470414 38898
rect 469794 2898 469826 3454
rect 470382 2898 470414 3454
rect 469794 -346 470414 2898
rect 469794 -902 469826 -346
rect 470382 -902 470414 -346
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690618 473546 691174
rect 474102 690618 474134 691174
rect 473514 655174 474134 690618
rect 473514 654618 473546 655174
rect 474102 654618 474134 655174
rect 473514 619174 474134 654618
rect 473514 618618 473546 619174
rect 474102 618618 474134 619174
rect 473514 583174 474134 618618
rect 473514 582618 473546 583174
rect 474102 582618 474134 583174
rect 473514 547174 474134 582618
rect 473514 546618 473546 547174
rect 474102 546618 474134 547174
rect 473514 511174 474134 546618
rect 473514 510618 473546 511174
rect 474102 510618 474134 511174
rect 473514 475174 474134 510618
rect 473514 474618 473546 475174
rect 474102 474618 474134 475174
rect 473514 439174 474134 474618
rect 473514 438618 473546 439174
rect 474102 438618 474134 439174
rect 473514 403174 474134 438618
rect 473514 402618 473546 403174
rect 474102 402618 474134 403174
rect 473514 367174 474134 402618
rect 473514 366618 473546 367174
rect 474102 366618 474134 367174
rect 473514 331174 474134 366618
rect 473514 330618 473546 331174
rect 474102 330618 474134 331174
rect 473514 295174 474134 330618
rect 473514 294618 473546 295174
rect 474102 294618 474134 295174
rect 473514 259174 474134 294618
rect 473514 258618 473546 259174
rect 474102 258618 474134 259174
rect 473514 223174 474134 258618
rect 473514 222618 473546 223174
rect 474102 222618 474134 223174
rect 473514 187174 474134 222618
rect 473514 186618 473546 187174
rect 474102 186618 474134 187174
rect 473514 151174 474134 186618
rect 473514 150618 473546 151174
rect 474102 150618 474134 151174
rect 473514 115174 474134 150618
rect 473514 114618 473546 115174
rect 474102 114618 474134 115174
rect 473514 79174 474134 114618
rect 473514 78618 473546 79174
rect 474102 78618 474134 79174
rect 473514 43174 474134 78618
rect 473514 42618 473546 43174
rect 474102 42618 474134 43174
rect 473514 7174 474134 42618
rect 473514 6618 473546 7174
rect 474102 6618 474134 7174
rect 473514 -2266 474134 6618
rect 473514 -2822 473546 -2266
rect 474102 -2822 474134 -2266
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694338 477266 694894
rect 477822 694338 477854 694894
rect 477234 658894 477854 694338
rect 477234 658338 477266 658894
rect 477822 658338 477854 658894
rect 477234 622894 477854 658338
rect 477234 622338 477266 622894
rect 477822 622338 477854 622894
rect 477234 586894 477854 622338
rect 477234 586338 477266 586894
rect 477822 586338 477854 586894
rect 477234 550894 477854 586338
rect 477234 550338 477266 550894
rect 477822 550338 477854 550894
rect 477234 514894 477854 550338
rect 477234 514338 477266 514894
rect 477822 514338 477854 514894
rect 477234 478894 477854 514338
rect 477234 478338 477266 478894
rect 477822 478338 477854 478894
rect 477234 442894 477854 478338
rect 477234 442338 477266 442894
rect 477822 442338 477854 442894
rect 477234 406894 477854 442338
rect 477234 406338 477266 406894
rect 477822 406338 477854 406894
rect 477234 370894 477854 406338
rect 477234 370338 477266 370894
rect 477822 370338 477854 370894
rect 477234 334894 477854 370338
rect 477234 334338 477266 334894
rect 477822 334338 477854 334894
rect 477234 298894 477854 334338
rect 477234 298338 477266 298894
rect 477822 298338 477854 298894
rect 477234 262894 477854 298338
rect 477234 262338 477266 262894
rect 477822 262338 477854 262894
rect 477234 226894 477854 262338
rect 477234 226338 477266 226894
rect 477822 226338 477854 226894
rect 477234 190894 477854 226338
rect 477234 190338 477266 190894
rect 477822 190338 477854 190894
rect 477234 154894 477854 190338
rect 477234 154338 477266 154894
rect 477822 154338 477854 154894
rect 477234 118894 477854 154338
rect 477234 118338 477266 118894
rect 477822 118338 477854 118894
rect 477234 82894 477854 118338
rect 477234 82338 477266 82894
rect 477822 82338 477854 82894
rect 477234 46894 477854 82338
rect 477234 46338 477266 46894
rect 477822 46338 477854 46894
rect 477234 10894 477854 46338
rect 477234 10338 477266 10894
rect 477822 10338 477854 10894
rect 477234 -4186 477854 10338
rect 477234 -4742 477266 -4186
rect 477822 -4742 477854 -4186
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711002 498986 711558
rect 499542 711002 499574 711558
rect 495234 709638 495854 709670
rect 495234 709082 495266 709638
rect 495822 709082 495854 709638
rect 491514 707718 492134 707750
rect 491514 707162 491546 707718
rect 492102 707162 492134 707718
rect 480954 698058 480986 698614
rect 481542 698058 481574 698614
rect 480954 662614 481574 698058
rect 480954 662058 480986 662614
rect 481542 662058 481574 662614
rect 480954 626614 481574 662058
rect 480954 626058 480986 626614
rect 481542 626058 481574 626614
rect 480954 590614 481574 626058
rect 480954 590058 480986 590614
rect 481542 590058 481574 590614
rect 480954 554614 481574 590058
rect 480954 554058 480986 554614
rect 481542 554058 481574 554614
rect 480954 518614 481574 554058
rect 480954 518058 480986 518614
rect 481542 518058 481574 518614
rect 480954 482614 481574 518058
rect 480954 482058 480986 482614
rect 481542 482058 481574 482614
rect 480954 446614 481574 482058
rect 480954 446058 480986 446614
rect 481542 446058 481574 446614
rect 480954 410614 481574 446058
rect 480954 410058 480986 410614
rect 481542 410058 481574 410614
rect 480954 374614 481574 410058
rect 480954 374058 480986 374614
rect 481542 374058 481574 374614
rect 480954 338614 481574 374058
rect 480954 338058 480986 338614
rect 481542 338058 481574 338614
rect 480954 302614 481574 338058
rect 480954 302058 480986 302614
rect 481542 302058 481574 302614
rect 480954 266614 481574 302058
rect 480954 266058 480986 266614
rect 481542 266058 481574 266614
rect 480954 230614 481574 266058
rect 480954 230058 480986 230614
rect 481542 230058 481574 230614
rect 480954 194614 481574 230058
rect 480954 194058 480986 194614
rect 481542 194058 481574 194614
rect 480954 158614 481574 194058
rect 480954 158058 480986 158614
rect 481542 158058 481574 158614
rect 480954 122614 481574 158058
rect 480954 122058 480986 122614
rect 481542 122058 481574 122614
rect 480954 86614 481574 122058
rect 480954 86058 480986 86614
rect 481542 86058 481574 86614
rect 480954 50614 481574 86058
rect 480954 50058 480986 50614
rect 481542 50058 481574 50614
rect 480954 14614 481574 50058
rect 480954 14058 480986 14614
rect 481542 14058 481574 14614
rect 462954 -7622 462986 -7066
rect 463542 -7622 463574 -7066
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705242 487826 705798
rect 488382 705242 488414 705798
rect 487794 669454 488414 705242
rect 487794 668898 487826 669454
rect 488382 668898 488414 669454
rect 487794 633454 488414 668898
rect 487794 632898 487826 633454
rect 488382 632898 488414 633454
rect 487794 597454 488414 632898
rect 487794 596898 487826 597454
rect 488382 596898 488414 597454
rect 487794 561454 488414 596898
rect 487794 560898 487826 561454
rect 488382 560898 488414 561454
rect 487794 525454 488414 560898
rect 487794 524898 487826 525454
rect 488382 524898 488414 525454
rect 487794 489454 488414 524898
rect 487794 488898 487826 489454
rect 488382 488898 488414 489454
rect 487794 453454 488414 488898
rect 487794 452898 487826 453454
rect 488382 452898 488414 453454
rect 487794 417454 488414 452898
rect 487794 416898 487826 417454
rect 488382 416898 488414 417454
rect 487794 381454 488414 416898
rect 487794 380898 487826 381454
rect 488382 380898 488414 381454
rect 487794 345454 488414 380898
rect 487794 344898 487826 345454
rect 488382 344898 488414 345454
rect 487794 309454 488414 344898
rect 487794 308898 487826 309454
rect 488382 308898 488414 309454
rect 487794 273454 488414 308898
rect 487794 272898 487826 273454
rect 488382 272898 488414 273454
rect 487794 237454 488414 272898
rect 487794 236898 487826 237454
rect 488382 236898 488414 237454
rect 487794 201454 488414 236898
rect 487794 200898 487826 201454
rect 488382 200898 488414 201454
rect 487794 165454 488414 200898
rect 487794 164898 487826 165454
rect 488382 164898 488414 165454
rect 487794 129454 488414 164898
rect 487794 128898 487826 129454
rect 488382 128898 488414 129454
rect 487794 93454 488414 128898
rect 487794 92898 487826 93454
rect 488382 92898 488414 93454
rect 487794 57454 488414 92898
rect 487794 56898 487826 57454
rect 488382 56898 488414 57454
rect 487794 21454 488414 56898
rect 487794 20898 487826 21454
rect 488382 20898 488414 21454
rect 487794 -1306 488414 20898
rect 487794 -1862 487826 -1306
rect 488382 -1862 488414 -1306
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672618 491546 673174
rect 492102 672618 492134 673174
rect 491514 637174 492134 672618
rect 491514 636618 491546 637174
rect 492102 636618 492134 637174
rect 491514 601174 492134 636618
rect 491514 600618 491546 601174
rect 492102 600618 492134 601174
rect 491514 565174 492134 600618
rect 491514 564618 491546 565174
rect 492102 564618 492134 565174
rect 491514 529174 492134 564618
rect 491514 528618 491546 529174
rect 492102 528618 492134 529174
rect 491514 493174 492134 528618
rect 491514 492618 491546 493174
rect 492102 492618 492134 493174
rect 491514 457174 492134 492618
rect 491514 456618 491546 457174
rect 492102 456618 492134 457174
rect 491514 421174 492134 456618
rect 491514 420618 491546 421174
rect 492102 420618 492134 421174
rect 491514 385174 492134 420618
rect 491514 384618 491546 385174
rect 492102 384618 492134 385174
rect 491514 349174 492134 384618
rect 491514 348618 491546 349174
rect 492102 348618 492134 349174
rect 491514 313174 492134 348618
rect 491514 312618 491546 313174
rect 492102 312618 492134 313174
rect 491514 277174 492134 312618
rect 491514 276618 491546 277174
rect 492102 276618 492134 277174
rect 491514 241174 492134 276618
rect 491514 240618 491546 241174
rect 492102 240618 492134 241174
rect 491514 205174 492134 240618
rect 491514 204618 491546 205174
rect 492102 204618 492134 205174
rect 491514 169174 492134 204618
rect 491514 168618 491546 169174
rect 492102 168618 492134 169174
rect 491514 133174 492134 168618
rect 491514 132618 491546 133174
rect 492102 132618 492134 133174
rect 491514 97174 492134 132618
rect 491514 96618 491546 97174
rect 492102 96618 492134 97174
rect 491514 61174 492134 96618
rect 491514 60618 491546 61174
rect 492102 60618 492134 61174
rect 491514 25174 492134 60618
rect 491514 24618 491546 25174
rect 492102 24618 492134 25174
rect 491514 -3226 492134 24618
rect 491514 -3782 491546 -3226
rect 492102 -3782 492134 -3226
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676338 495266 676894
rect 495822 676338 495854 676894
rect 495234 640894 495854 676338
rect 495234 640338 495266 640894
rect 495822 640338 495854 640894
rect 495234 604894 495854 640338
rect 495234 604338 495266 604894
rect 495822 604338 495854 604894
rect 495234 568894 495854 604338
rect 495234 568338 495266 568894
rect 495822 568338 495854 568894
rect 495234 532894 495854 568338
rect 495234 532338 495266 532894
rect 495822 532338 495854 532894
rect 495234 496894 495854 532338
rect 495234 496338 495266 496894
rect 495822 496338 495854 496894
rect 495234 460894 495854 496338
rect 495234 460338 495266 460894
rect 495822 460338 495854 460894
rect 495234 424894 495854 460338
rect 495234 424338 495266 424894
rect 495822 424338 495854 424894
rect 495234 388894 495854 424338
rect 495234 388338 495266 388894
rect 495822 388338 495854 388894
rect 495234 352894 495854 388338
rect 495234 352338 495266 352894
rect 495822 352338 495854 352894
rect 495234 316894 495854 352338
rect 495234 316338 495266 316894
rect 495822 316338 495854 316894
rect 495234 280894 495854 316338
rect 495234 280338 495266 280894
rect 495822 280338 495854 280894
rect 495234 244894 495854 280338
rect 495234 244338 495266 244894
rect 495822 244338 495854 244894
rect 495234 208894 495854 244338
rect 495234 208338 495266 208894
rect 495822 208338 495854 208894
rect 495234 172894 495854 208338
rect 495234 172338 495266 172894
rect 495822 172338 495854 172894
rect 495234 136894 495854 172338
rect 495234 136338 495266 136894
rect 495822 136338 495854 136894
rect 495234 100894 495854 136338
rect 495234 100338 495266 100894
rect 495822 100338 495854 100894
rect 495234 64894 495854 100338
rect 495234 64338 495266 64894
rect 495822 64338 495854 64894
rect 495234 28894 495854 64338
rect 495234 28338 495266 28894
rect 495822 28338 495854 28894
rect 495234 -5146 495854 28338
rect 495234 -5702 495266 -5146
rect 495822 -5702 495854 -5146
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710042 516986 710598
rect 517542 710042 517574 710598
rect 513234 708678 513854 709670
rect 513234 708122 513266 708678
rect 513822 708122 513854 708678
rect 509514 706758 510134 707750
rect 509514 706202 509546 706758
rect 510102 706202 510134 706758
rect 498954 680058 498986 680614
rect 499542 680058 499574 680614
rect 498954 644614 499574 680058
rect 498954 644058 498986 644614
rect 499542 644058 499574 644614
rect 498954 608614 499574 644058
rect 498954 608058 498986 608614
rect 499542 608058 499574 608614
rect 498954 572614 499574 608058
rect 498954 572058 498986 572614
rect 499542 572058 499574 572614
rect 498954 536614 499574 572058
rect 498954 536058 498986 536614
rect 499542 536058 499574 536614
rect 498954 500614 499574 536058
rect 498954 500058 498986 500614
rect 499542 500058 499574 500614
rect 498954 464614 499574 500058
rect 498954 464058 498986 464614
rect 499542 464058 499574 464614
rect 498954 428614 499574 464058
rect 498954 428058 498986 428614
rect 499542 428058 499574 428614
rect 498954 392614 499574 428058
rect 498954 392058 498986 392614
rect 499542 392058 499574 392614
rect 498954 356614 499574 392058
rect 498954 356058 498986 356614
rect 499542 356058 499574 356614
rect 498954 320614 499574 356058
rect 498954 320058 498986 320614
rect 499542 320058 499574 320614
rect 498954 284614 499574 320058
rect 498954 284058 498986 284614
rect 499542 284058 499574 284614
rect 498954 248614 499574 284058
rect 498954 248058 498986 248614
rect 499542 248058 499574 248614
rect 498954 212614 499574 248058
rect 498954 212058 498986 212614
rect 499542 212058 499574 212614
rect 498954 176614 499574 212058
rect 498954 176058 498986 176614
rect 499542 176058 499574 176614
rect 498954 140614 499574 176058
rect 498954 140058 498986 140614
rect 499542 140058 499574 140614
rect 498954 104614 499574 140058
rect 498954 104058 498986 104614
rect 499542 104058 499574 104614
rect 498954 68614 499574 104058
rect 498954 68058 498986 68614
rect 499542 68058 499574 68614
rect 498954 32614 499574 68058
rect 498954 32058 498986 32614
rect 499542 32058 499574 32614
rect 480954 -6662 480986 -6106
rect 481542 -6662 481574 -6106
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704282 505826 704838
rect 506382 704282 506414 704838
rect 505794 687454 506414 704282
rect 505794 686898 505826 687454
rect 506382 686898 506414 687454
rect 505794 651454 506414 686898
rect 505794 650898 505826 651454
rect 506382 650898 506414 651454
rect 505794 615454 506414 650898
rect 505794 614898 505826 615454
rect 506382 614898 506414 615454
rect 505794 579454 506414 614898
rect 505794 578898 505826 579454
rect 506382 578898 506414 579454
rect 505794 543454 506414 578898
rect 505794 542898 505826 543454
rect 506382 542898 506414 543454
rect 505794 507454 506414 542898
rect 505794 506898 505826 507454
rect 506382 506898 506414 507454
rect 505794 471454 506414 506898
rect 505794 470898 505826 471454
rect 506382 470898 506414 471454
rect 505794 435454 506414 470898
rect 505794 434898 505826 435454
rect 506382 434898 506414 435454
rect 505794 399454 506414 434898
rect 505794 398898 505826 399454
rect 506382 398898 506414 399454
rect 505794 363454 506414 398898
rect 505794 362898 505826 363454
rect 506382 362898 506414 363454
rect 505794 327454 506414 362898
rect 505794 326898 505826 327454
rect 506382 326898 506414 327454
rect 505794 291454 506414 326898
rect 505794 290898 505826 291454
rect 506382 290898 506414 291454
rect 505794 255454 506414 290898
rect 505794 254898 505826 255454
rect 506382 254898 506414 255454
rect 505794 219454 506414 254898
rect 505794 218898 505826 219454
rect 506382 218898 506414 219454
rect 505794 183454 506414 218898
rect 505794 182898 505826 183454
rect 506382 182898 506414 183454
rect 505794 147454 506414 182898
rect 505794 146898 505826 147454
rect 506382 146898 506414 147454
rect 505794 111454 506414 146898
rect 505794 110898 505826 111454
rect 506382 110898 506414 111454
rect 505794 75454 506414 110898
rect 505794 74898 505826 75454
rect 506382 74898 506414 75454
rect 505794 39454 506414 74898
rect 505794 38898 505826 39454
rect 506382 38898 506414 39454
rect 505794 3454 506414 38898
rect 505794 2898 505826 3454
rect 506382 2898 506414 3454
rect 505794 -346 506414 2898
rect 505794 -902 505826 -346
rect 506382 -902 506414 -346
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690618 509546 691174
rect 510102 690618 510134 691174
rect 509514 655174 510134 690618
rect 509514 654618 509546 655174
rect 510102 654618 510134 655174
rect 509514 619174 510134 654618
rect 509514 618618 509546 619174
rect 510102 618618 510134 619174
rect 509514 583174 510134 618618
rect 509514 582618 509546 583174
rect 510102 582618 510134 583174
rect 509514 547174 510134 582618
rect 509514 546618 509546 547174
rect 510102 546618 510134 547174
rect 509514 511174 510134 546618
rect 509514 510618 509546 511174
rect 510102 510618 510134 511174
rect 509514 475174 510134 510618
rect 509514 474618 509546 475174
rect 510102 474618 510134 475174
rect 509514 439174 510134 474618
rect 509514 438618 509546 439174
rect 510102 438618 510134 439174
rect 509514 403174 510134 438618
rect 509514 402618 509546 403174
rect 510102 402618 510134 403174
rect 509514 367174 510134 402618
rect 509514 366618 509546 367174
rect 510102 366618 510134 367174
rect 509514 331174 510134 366618
rect 509514 330618 509546 331174
rect 510102 330618 510134 331174
rect 509514 295174 510134 330618
rect 509514 294618 509546 295174
rect 510102 294618 510134 295174
rect 509514 259174 510134 294618
rect 509514 258618 509546 259174
rect 510102 258618 510134 259174
rect 509514 223174 510134 258618
rect 509514 222618 509546 223174
rect 510102 222618 510134 223174
rect 509514 187174 510134 222618
rect 509514 186618 509546 187174
rect 510102 186618 510134 187174
rect 509514 151174 510134 186618
rect 509514 150618 509546 151174
rect 510102 150618 510134 151174
rect 509514 115174 510134 150618
rect 509514 114618 509546 115174
rect 510102 114618 510134 115174
rect 509514 79174 510134 114618
rect 509514 78618 509546 79174
rect 510102 78618 510134 79174
rect 509514 43174 510134 78618
rect 509514 42618 509546 43174
rect 510102 42618 510134 43174
rect 509514 7174 510134 42618
rect 509514 6618 509546 7174
rect 510102 6618 510134 7174
rect 509514 -2266 510134 6618
rect 509514 -2822 509546 -2266
rect 510102 -2822 510134 -2266
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694338 513266 694894
rect 513822 694338 513854 694894
rect 513234 658894 513854 694338
rect 513234 658338 513266 658894
rect 513822 658338 513854 658894
rect 513234 622894 513854 658338
rect 513234 622338 513266 622894
rect 513822 622338 513854 622894
rect 513234 586894 513854 622338
rect 513234 586338 513266 586894
rect 513822 586338 513854 586894
rect 513234 550894 513854 586338
rect 513234 550338 513266 550894
rect 513822 550338 513854 550894
rect 513234 514894 513854 550338
rect 513234 514338 513266 514894
rect 513822 514338 513854 514894
rect 513234 478894 513854 514338
rect 513234 478338 513266 478894
rect 513822 478338 513854 478894
rect 513234 442894 513854 478338
rect 513234 442338 513266 442894
rect 513822 442338 513854 442894
rect 513234 406894 513854 442338
rect 513234 406338 513266 406894
rect 513822 406338 513854 406894
rect 513234 370894 513854 406338
rect 513234 370338 513266 370894
rect 513822 370338 513854 370894
rect 513234 334894 513854 370338
rect 513234 334338 513266 334894
rect 513822 334338 513854 334894
rect 513234 298894 513854 334338
rect 513234 298338 513266 298894
rect 513822 298338 513854 298894
rect 513234 262894 513854 298338
rect 513234 262338 513266 262894
rect 513822 262338 513854 262894
rect 513234 226894 513854 262338
rect 513234 226338 513266 226894
rect 513822 226338 513854 226894
rect 513234 190894 513854 226338
rect 513234 190338 513266 190894
rect 513822 190338 513854 190894
rect 513234 154894 513854 190338
rect 513234 154338 513266 154894
rect 513822 154338 513854 154894
rect 513234 118894 513854 154338
rect 513234 118338 513266 118894
rect 513822 118338 513854 118894
rect 513234 82894 513854 118338
rect 513234 82338 513266 82894
rect 513822 82338 513854 82894
rect 513234 46894 513854 82338
rect 513234 46338 513266 46894
rect 513822 46338 513854 46894
rect 513234 10894 513854 46338
rect 513234 10338 513266 10894
rect 513822 10338 513854 10894
rect 513234 -4186 513854 10338
rect 513234 -4742 513266 -4186
rect 513822 -4742 513854 -4186
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711002 534986 711558
rect 535542 711002 535574 711558
rect 531234 709638 531854 709670
rect 531234 709082 531266 709638
rect 531822 709082 531854 709638
rect 527514 707718 528134 707750
rect 527514 707162 527546 707718
rect 528102 707162 528134 707718
rect 516954 698058 516986 698614
rect 517542 698058 517574 698614
rect 516954 662614 517574 698058
rect 516954 662058 516986 662614
rect 517542 662058 517574 662614
rect 516954 626614 517574 662058
rect 516954 626058 516986 626614
rect 517542 626058 517574 626614
rect 516954 590614 517574 626058
rect 516954 590058 516986 590614
rect 517542 590058 517574 590614
rect 516954 554614 517574 590058
rect 516954 554058 516986 554614
rect 517542 554058 517574 554614
rect 516954 518614 517574 554058
rect 516954 518058 516986 518614
rect 517542 518058 517574 518614
rect 516954 482614 517574 518058
rect 516954 482058 516986 482614
rect 517542 482058 517574 482614
rect 516954 446614 517574 482058
rect 516954 446058 516986 446614
rect 517542 446058 517574 446614
rect 516954 410614 517574 446058
rect 516954 410058 516986 410614
rect 517542 410058 517574 410614
rect 516954 374614 517574 410058
rect 516954 374058 516986 374614
rect 517542 374058 517574 374614
rect 516954 338614 517574 374058
rect 516954 338058 516986 338614
rect 517542 338058 517574 338614
rect 516954 302614 517574 338058
rect 516954 302058 516986 302614
rect 517542 302058 517574 302614
rect 516954 266614 517574 302058
rect 516954 266058 516986 266614
rect 517542 266058 517574 266614
rect 516954 230614 517574 266058
rect 516954 230058 516986 230614
rect 517542 230058 517574 230614
rect 516954 194614 517574 230058
rect 516954 194058 516986 194614
rect 517542 194058 517574 194614
rect 516954 158614 517574 194058
rect 516954 158058 516986 158614
rect 517542 158058 517574 158614
rect 516954 122614 517574 158058
rect 516954 122058 516986 122614
rect 517542 122058 517574 122614
rect 516954 86614 517574 122058
rect 516954 86058 516986 86614
rect 517542 86058 517574 86614
rect 516954 50614 517574 86058
rect 516954 50058 516986 50614
rect 517542 50058 517574 50614
rect 516954 14614 517574 50058
rect 516954 14058 516986 14614
rect 517542 14058 517574 14614
rect 498954 -7622 498986 -7066
rect 499542 -7622 499574 -7066
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705242 523826 705798
rect 524382 705242 524414 705798
rect 523794 669454 524414 705242
rect 523794 668898 523826 669454
rect 524382 668898 524414 669454
rect 523794 633454 524414 668898
rect 523794 632898 523826 633454
rect 524382 632898 524414 633454
rect 523794 597454 524414 632898
rect 523794 596898 523826 597454
rect 524382 596898 524414 597454
rect 523794 561454 524414 596898
rect 523794 560898 523826 561454
rect 524382 560898 524414 561454
rect 523794 525454 524414 560898
rect 523794 524898 523826 525454
rect 524382 524898 524414 525454
rect 523794 489454 524414 524898
rect 523794 488898 523826 489454
rect 524382 488898 524414 489454
rect 523794 453454 524414 488898
rect 523794 452898 523826 453454
rect 524382 452898 524414 453454
rect 523794 417454 524414 452898
rect 523794 416898 523826 417454
rect 524382 416898 524414 417454
rect 523794 381454 524414 416898
rect 523794 380898 523826 381454
rect 524382 380898 524414 381454
rect 523794 345454 524414 380898
rect 523794 344898 523826 345454
rect 524382 344898 524414 345454
rect 523794 309454 524414 344898
rect 523794 308898 523826 309454
rect 524382 308898 524414 309454
rect 523794 273454 524414 308898
rect 523794 272898 523826 273454
rect 524382 272898 524414 273454
rect 523794 237454 524414 272898
rect 523794 236898 523826 237454
rect 524382 236898 524414 237454
rect 523794 201454 524414 236898
rect 523794 200898 523826 201454
rect 524382 200898 524414 201454
rect 523794 165454 524414 200898
rect 523794 164898 523826 165454
rect 524382 164898 524414 165454
rect 523794 129454 524414 164898
rect 523794 128898 523826 129454
rect 524382 128898 524414 129454
rect 523794 93454 524414 128898
rect 523794 92898 523826 93454
rect 524382 92898 524414 93454
rect 523794 57454 524414 92898
rect 523794 56898 523826 57454
rect 524382 56898 524414 57454
rect 523794 21454 524414 56898
rect 523794 20898 523826 21454
rect 524382 20898 524414 21454
rect 523794 -1306 524414 20898
rect 523794 -1862 523826 -1306
rect 524382 -1862 524414 -1306
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672618 527546 673174
rect 528102 672618 528134 673174
rect 527514 637174 528134 672618
rect 527514 636618 527546 637174
rect 528102 636618 528134 637174
rect 527514 601174 528134 636618
rect 527514 600618 527546 601174
rect 528102 600618 528134 601174
rect 527514 565174 528134 600618
rect 527514 564618 527546 565174
rect 528102 564618 528134 565174
rect 527514 529174 528134 564618
rect 527514 528618 527546 529174
rect 528102 528618 528134 529174
rect 527514 493174 528134 528618
rect 527514 492618 527546 493174
rect 528102 492618 528134 493174
rect 527514 457174 528134 492618
rect 527514 456618 527546 457174
rect 528102 456618 528134 457174
rect 527514 421174 528134 456618
rect 527514 420618 527546 421174
rect 528102 420618 528134 421174
rect 527514 385174 528134 420618
rect 527514 384618 527546 385174
rect 528102 384618 528134 385174
rect 527514 349174 528134 384618
rect 527514 348618 527546 349174
rect 528102 348618 528134 349174
rect 527514 313174 528134 348618
rect 527514 312618 527546 313174
rect 528102 312618 528134 313174
rect 527514 277174 528134 312618
rect 527514 276618 527546 277174
rect 528102 276618 528134 277174
rect 527514 241174 528134 276618
rect 527514 240618 527546 241174
rect 528102 240618 528134 241174
rect 527514 205174 528134 240618
rect 527514 204618 527546 205174
rect 528102 204618 528134 205174
rect 527514 169174 528134 204618
rect 527514 168618 527546 169174
rect 528102 168618 528134 169174
rect 527514 133174 528134 168618
rect 527514 132618 527546 133174
rect 528102 132618 528134 133174
rect 527514 97174 528134 132618
rect 527514 96618 527546 97174
rect 528102 96618 528134 97174
rect 527514 61174 528134 96618
rect 527514 60618 527546 61174
rect 528102 60618 528134 61174
rect 527514 25174 528134 60618
rect 527514 24618 527546 25174
rect 528102 24618 528134 25174
rect 527514 -3226 528134 24618
rect 527514 -3782 527546 -3226
rect 528102 -3782 528134 -3226
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676338 531266 676894
rect 531822 676338 531854 676894
rect 531234 640894 531854 676338
rect 531234 640338 531266 640894
rect 531822 640338 531854 640894
rect 531234 604894 531854 640338
rect 531234 604338 531266 604894
rect 531822 604338 531854 604894
rect 531234 568894 531854 604338
rect 531234 568338 531266 568894
rect 531822 568338 531854 568894
rect 531234 532894 531854 568338
rect 531234 532338 531266 532894
rect 531822 532338 531854 532894
rect 531234 496894 531854 532338
rect 531234 496338 531266 496894
rect 531822 496338 531854 496894
rect 531234 460894 531854 496338
rect 531234 460338 531266 460894
rect 531822 460338 531854 460894
rect 531234 424894 531854 460338
rect 531234 424338 531266 424894
rect 531822 424338 531854 424894
rect 531234 388894 531854 424338
rect 531234 388338 531266 388894
rect 531822 388338 531854 388894
rect 531234 352894 531854 388338
rect 531234 352338 531266 352894
rect 531822 352338 531854 352894
rect 531234 316894 531854 352338
rect 531234 316338 531266 316894
rect 531822 316338 531854 316894
rect 531234 280894 531854 316338
rect 531234 280338 531266 280894
rect 531822 280338 531854 280894
rect 531234 244894 531854 280338
rect 531234 244338 531266 244894
rect 531822 244338 531854 244894
rect 531234 208894 531854 244338
rect 531234 208338 531266 208894
rect 531822 208338 531854 208894
rect 531234 172894 531854 208338
rect 531234 172338 531266 172894
rect 531822 172338 531854 172894
rect 531234 136894 531854 172338
rect 531234 136338 531266 136894
rect 531822 136338 531854 136894
rect 531234 100894 531854 136338
rect 531234 100338 531266 100894
rect 531822 100338 531854 100894
rect 531234 64894 531854 100338
rect 531234 64338 531266 64894
rect 531822 64338 531854 64894
rect 531234 28894 531854 64338
rect 531234 28338 531266 28894
rect 531822 28338 531854 28894
rect 531234 -5146 531854 28338
rect 531234 -5702 531266 -5146
rect 531822 -5702 531854 -5146
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710042 552986 710598
rect 553542 710042 553574 710598
rect 549234 708678 549854 709670
rect 549234 708122 549266 708678
rect 549822 708122 549854 708678
rect 545514 706758 546134 707750
rect 545514 706202 545546 706758
rect 546102 706202 546134 706758
rect 534954 680058 534986 680614
rect 535542 680058 535574 680614
rect 534954 644614 535574 680058
rect 534954 644058 534986 644614
rect 535542 644058 535574 644614
rect 534954 608614 535574 644058
rect 534954 608058 534986 608614
rect 535542 608058 535574 608614
rect 534954 572614 535574 608058
rect 534954 572058 534986 572614
rect 535542 572058 535574 572614
rect 534954 536614 535574 572058
rect 534954 536058 534986 536614
rect 535542 536058 535574 536614
rect 534954 500614 535574 536058
rect 534954 500058 534986 500614
rect 535542 500058 535574 500614
rect 534954 464614 535574 500058
rect 534954 464058 534986 464614
rect 535542 464058 535574 464614
rect 534954 428614 535574 464058
rect 534954 428058 534986 428614
rect 535542 428058 535574 428614
rect 534954 392614 535574 428058
rect 534954 392058 534986 392614
rect 535542 392058 535574 392614
rect 534954 356614 535574 392058
rect 534954 356058 534986 356614
rect 535542 356058 535574 356614
rect 534954 320614 535574 356058
rect 534954 320058 534986 320614
rect 535542 320058 535574 320614
rect 534954 284614 535574 320058
rect 534954 284058 534986 284614
rect 535542 284058 535574 284614
rect 534954 248614 535574 284058
rect 534954 248058 534986 248614
rect 535542 248058 535574 248614
rect 534954 212614 535574 248058
rect 534954 212058 534986 212614
rect 535542 212058 535574 212614
rect 534954 176614 535574 212058
rect 534954 176058 534986 176614
rect 535542 176058 535574 176614
rect 534954 140614 535574 176058
rect 534954 140058 534986 140614
rect 535542 140058 535574 140614
rect 534954 104614 535574 140058
rect 534954 104058 534986 104614
rect 535542 104058 535574 104614
rect 534954 68614 535574 104058
rect 534954 68058 534986 68614
rect 535542 68058 535574 68614
rect 534954 32614 535574 68058
rect 534954 32058 534986 32614
rect 535542 32058 535574 32614
rect 516954 -6662 516986 -6106
rect 517542 -6662 517574 -6106
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704282 541826 704838
rect 542382 704282 542414 704838
rect 541794 687454 542414 704282
rect 541794 686898 541826 687454
rect 542382 686898 542414 687454
rect 541794 651454 542414 686898
rect 541794 650898 541826 651454
rect 542382 650898 542414 651454
rect 541794 615454 542414 650898
rect 541794 614898 541826 615454
rect 542382 614898 542414 615454
rect 541794 579454 542414 614898
rect 541794 578898 541826 579454
rect 542382 578898 542414 579454
rect 541794 543454 542414 578898
rect 541794 542898 541826 543454
rect 542382 542898 542414 543454
rect 541794 507454 542414 542898
rect 541794 506898 541826 507454
rect 542382 506898 542414 507454
rect 541794 471454 542414 506898
rect 541794 470898 541826 471454
rect 542382 470898 542414 471454
rect 541794 435454 542414 470898
rect 541794 434898 541826 435454
rect 542382 434898 542414 435454
rect 541794 399454 542414 434898
rect 541794 398898 541826 399454
rect 542382 398898 542414 399454
rect 541794 363454 542414 398898
rect 541794 362898 541826 363454
rect 542382 362898 542414 363454
rect 541794 327454 542414 362898
rect 541794 326898 541826 327454
rect 542382 326898 542414 327454
rect 541794 291454 542414 326898
rect 541794 290898 541826 291454
rect 542382 290898 542414 291454
rect 541794 255454 542414 290898
rect 541794 254898 541826 255454
rect 542382 254898 542414 255454
rect 541794 219454 542414 254898
rect 541794 218898 541826 219454
rect 542382 218898 542414 219454
rect 541794 183454 542414 218898
rect 541794 182898 541826 183454
rect 542382 182898 542414 183454
rect 541794 147454 542414 182898
rect 541794 146898 541826 147454
rect 542382 146898 542414 147454
rect 541794 111454 542414 146898
rect 541794 110898 541826 111454
rect 542382 110898 542414 111454
rect 541794 75454 542414 110898
rect 541794 74898 541826 75454
rect 542382 74898 542414 75454
rect 541794 39454 542414 74898
rect 541794 38898 541826 39454
rect 542382 38898 542414 39454
rect 541794 3454 542414 38898
rect 541794 2898 541826 3454
rect 542382 2898 542414 3454
rect 541794 -346 542414 2898
rect 541794 -902 541826 -346
rect 542382 -902 542414 -346
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690618 545546 691174
rect 546102 690618 546134 691174
rect 545514 655174 546134 690618
rect 545514 654618 545546 655174
rect 546102 654618 546134 655174
rect 545514 619174 546134 654618
rect 545514 618618 545546 619174
rect 546102 618618 546134 619174
rect 545514 583174 546134 618618
rect 545514 582618 545546 583174
rect 546102 582618 546134 583174
rect 545514 547174 546134 582618
rect 545514 546618 545546 547174
rect 546102 546618 546134 547174
rect 545514 511174 546134 546618
rect 545514 510618 545546 511174
rect 546102 510618 546134 511174
rect 545514 475174 546134 510618
rect 545514 474618 545546 475174
rect 546102 474618 546134 475174
rect 545514 439174 546134 474618
rect 545514 438618 545546 439174
rect 546102 438618 546134 439174
rect 545514 403174 546134 438618
rect 545514 402618 545546 403174
rect 546102 402618 546134 403174
rect 545514 367174 546134 402618
rect 545514 366618 545546 367174
rect 546102 366618 546134 367174
rect 545514 331174 546134 366618
rect 545514 330618 545546 331174
rect 546102 330618 546134 331174
rect 545514 295174 546134 330618
rect 545514 294618 545546 295174
rect 546102 294618 546134 295174
rect 545514 259174 546134 294618
rect 545514 258618 545546 259174
rect 546102 258618 546134 259174
rect 545514 223174 546134 258618
rect 545514 222618 545546 223174
rect 546102 222618 546134 223174
rect 545514 187174 546134 222618
rect 545514 186618 545546 187174
rect 546102 186618 546134 187174
rect 545514 151174 546134 186618
rect 545514 150618 545546 151174
rect 546102 150618 546134 151174
rect 545514 115174 546134 150618
rect 545514 114618 545546 115174
rect 546102 114618 546134 115174
rect 545514 79174 546134 114618
rect 545514 78618 545546 79174
rect 546102 78618 546134 79174
rect 545514 43174 546134 78618
rect 545514 42618 545546 43174
rect 546102 42618 546134 43174
rect 545514 7174 546134 42618
rect 545514 6618 545546 7174
rect 546102 6618 546134 7174
rect 545514 -2266 546134 6618
rect 545514 -2822 545546 -2266
rect 546102 -2822 546134 -2266
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694338 549266 694894
rect 549822 694338 549854 694894
rect 549234 658894 549854 694338
rect 549234 658338 549266 658894
rect 549822 658338 549854 658894
rect 549234 622894 549854 658338
rect 549234 622338 549266 622894
rect 549822 622338 549854 622894
rect 549234 586894 549854 622338
rect 549234 586338 549266 586894
rect 549822 586338 549854 586894
rect 549234 550894 549854 586338
rect 549234 550338 549266 550894
rect 549822 550338 549854 550894
rect 549234 514894 549854 550338
rect 549234 514338 549266 514894
rect 549822 514338 549854 514894
rect 549234 478894 549854 514338
rect 549234 478338 549266 478894
rect 549822 478338 549854 478894
rect 549234 442894 549854 478338
rect 549234 442338 549266 442894
rect 549822 442338 549854 442894
rect 549234 406894 549854 442338
rect 549234 406338 549266 406894
rect 549822 406338 549854 406894
rect 549234 370894 549854 406338
rect 549234 370338 549266 370894
rect 549822 370338 549854 370894
rect 549234 334894 549854 370338
rect 549234 334338 549266 334894
rect 549822 334338 549854 334894
rect 549234 298894 549854 334338
rect 549234 298338 549266 298894
rect 549822 298338 549854 298894
rect 549234 262894 549854 298338
rect 549234 262338 549266 262894
rect 549822 262338 549854 262894
rect 549234 226894 549854 262338
rect 549234 226338 549266 226894
rect 549822 226338 549854 226894
rect 549234 190894 549854 226338
rect 549234 190338 549266 190894
rect 549822 190338 549854 190894
rect 549234 154894 549854 190338
rect 549234 154338 549266 154894
rect 549822 154338 549854 154894
rect 549234 118894 549854 154338
rect 549234 118338 549266 118894
rect 549822 118338 549854 118894
rect 549234 82894 549854 118338
rect 549234 82338 549266 82894
rect 549822 82338 549854 82894
rect 549234 46894 549854 82338
rect 549234 46338 549266 46894
rect 549822 46338 549854 46894
rect 549234 10894 549854 46338
rect 549234 10338 549266 10894
rect 549822 10338 549854 10894
rect 549234 -4186 549854 10338
rect 549234 -4742 549266 -4186
rect 549822 -4742 549854 -4186
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711002 570986 711558
rect 571542 711002 571574 711558
rect 567234 709638 567854 709670
rect 567234 709082 567266 709638
rect 567822 709082 567854 709638
rect 563514 707718 564134 707750
rect 563514 707162 563546 707718
rect 564102 707162 564134 707718
rect 552954 698058 552986 698614
rect 553542 698058 553574 698614
rect 552954 662614 553574 698058
rect 552954 662058 552986 662614
rect 553542 662058 553574 662614
rect 552954 626614 553574 662058
rect 552954 626058 552986 626614
rect 553542 626058 553574 626614
rect 552954 590614 553574 626058
rect 552954 590058 552986 590614
rect 553542 590058 553574 590614
rect 552954 554614 553574 590058
rect 552954 554058 552986 554614
rect 553542 554058 553574 554614
rect 552954 518614 553574 554058
rect 552954 518058 552986 518614
rect 553542 518058 553574 518614
rect 552954 482614 553574 518058
rect 552954 482058 552986 482614
rect 553542 482058 553574 482614
rect 552954 446614 553574 482058
rect 552954 446058 552986 446614
rect 553542 446058 553574 446614
rect 552954 410614 553574 446058
rect 552954 410058 552986 410614
rect 553542 410058 553574 410614
rect 552954 374614 553574 410058
rect 552954 374058 552986 374614
rect 553542 374058 553574 374614
rect 552954 338614 553574 374058
rect 552954 338058 552986 338614
rect 553542 338058 553574 338614
rect 552954 302614 553574 338058
rect 552954 302058 552986 302614
rect 553542 302058 553574 302614
rect 552954 266614 553574 302058
rect 552954 266058 552986 266614
rect 553542 266058 553574 266614
rect 552954 230614 553574 266058
rect 552954 230058 552986 230614
rect 553542 230058 553574 230614
rect 552954 194614 553574 230058
rect 552954 194058 552986 194614
rect 553542 194058 553574 194614
rect 552954 158614 553574 194058
rect 552954 158058 552986 158614
rect 553542 158058 553574 158614
rect 552954 122614 553574 158058
rect 552954 122058 552986 122614
rect 553542 122058 553574 122614
rect 552954 86614 553574 122058
rect 552954 86058 552986 86614
rect 553542 86058 553574 86614
rect 552954 50614 553574 86058
rect 552954 50058 552986 50614
rect 553542 50058 553574 50614
rect 552954 14614 553574 50058
rect 552954 14058 552986 14614
rect 553542 14058 553574 14614
rect 534954 -7622 534986 -7066
rect 535542 -7622 535574 -7066
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705242 559826 705798
rect 560382 705242 560414 705798
rect 559794 669454 560414 705242
rect 559794 668898 559826 669454
rect 560382 668898 560414 669454
rect 559794 633454 560414 668898
rect 559794 632898 559826 633454
rect 560382 632898 560414 633454
rect 559794 597454 560414 632898
rect 559794 596898 559826 597454
rect 560382 596898 560414 597454
rect 559794 561454 560414 596898
rect 559794 560898 559826 561454
rect 560382 560898 560414 561454
rect 559794 525454 560414 560898
rect 559794 524898 559826 525454
rect 560382 524898 560414 525454
rect 559794 489454 560414 524898
rect 559794 488898 559826 489454
rect 560382 488898 560414 489454
rect 559794 453454 560414 488898
rect 559794 452898 559826 453454
rect 560382 452898 560414 453454
rect 559794 417454 560414 452898
rect 559794 416898 559826 417454
rect 560382 416898 560414 417454
rect 559794 381454 560414 416898
rect 559794 380898 559826 381454
rect 560382 380898 560414 381454
rect 559794 345454 560414 380898
rect 559794 344898 559826 345454
rect 560382 344898 560414 345454
rect 559794 309454 560414 344898
rect 559794 308898 559826 309454
rect 560382 308898 560414 309454
rect 559794 273454 560414 308898
rect 559794 272898 559826 273454
rect 560382 272898 560414 273454
rect 559794 237454 560414 272898
rect 559794 236898 559826 237454
rect 560382 236898 560414 237454
rect 559794 201454 560414 236898
rect 559794 200898 559826 201454
rect 560382 200898 560414 201454
rect 559794 165454 560414 200898
rect 559794 164898 559826 165454
rect 560382 164898 560414 165454
rect 559794 129454 560414 164898
rect 559794 128898 559826 129454
rect 560382 128898 560414 129454
rect 559794 93454 560414 128898
rect 559794 92898 559826 93454
rect 560382 92898 560414 93454
rect 559794 57454 560414 92898
rect 559794 56898 559826 57454
rect 560382 56898 560414 57454
rect 559794 21454 560414 56898
rect 559794 20898 559826 21454
rect 560382 20898 560414 21454
rect 559794 -1306 560414 20898
rect 559794 -1862 559826 -1306
rect 560382 -1862 560414 -1306
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672618 563546 673174
rect 564102 672618 564134 673174
rect 563514 637174 564134 672618
rect 563514 636618 563546 637174
rect 564102 636618 564134 637174
rect 563514 601174 564134 636618
rect 563514 600618 563546 601174
rect 564102 600618 564134 601174
rect 563514 565174 564134 600618
rect 563514 564618 563546 565174
rect 564102 564618 564134 565174
rect 563514 529174 564134 564618
rect 563514 528618 563546 529174
rect 564102 528618 564134 529174
rect 563514 493174 564134 528618
rect 563514 492618 563546 493174
rect 564102 492618 564134 493174
rect 563514 457174 564134 492618
rect 563514 456618 563546 457174
rect 564102 456618 564134 457174
rect 563514 421174 564134 456618
rect 563514 420618 563546 421174
rect 564102 420618 564134 421174
rect 563514 385174 564134 420618
rect 563514 384618 563546 385174
rect 564102 384618 564134 385174
rect 563514 349174 564134 384618
rect 563514 348618 563546 349174
rect 564102 348618 564134 349174
rect 563514 313174 564134 348618
rect 563514 312618 563546 313174
rect 564102 312618 564134 313174
rect 563514 277174 564134 312618
rect 563514 276618 563546 277174
rect 564102 276618 564134 277174
rect 563514 241174 564134 276618
rect 563514 240618 563546 241174
rect 564102 240618 564134 241174
rect 563514 205174 564134 240618
rect 563514 204618 563546 205174
rect 564102 204618 564134 205174
rect 563514 169174 564134 204618
rect 563514 168618 563546 169174
rect 564102 168618 564134 169174
rect 563514 133174 564134 168618
rect 563514 132618 563546 133174
rect 564102 132618 564134 133174
rect 563514 97174 564134 132618
rect 563514 96618 563546 97174
rect 564102 96618 564134 97174
rect 563514 61174 564134 96618
rect 563514 60618 563546 61174
rect 564102 60618 564134 61174
rect 563514 25174 564134 60618
rect 563514 24618 563546 25174
rect 564102 24618 564134 25174
rect 563514 -3226 564134 24618
rect 563514 -3782 563546 -3226
rect 564102 -3782 564134 -3226
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676338 567266 676894
rect 567822 676338 567854 676894
rect 567234 640894 567854 676338
rect 567234 640338 567266 640894
rect 567822 640338 567854 640894
rect 567234 604894 567854 640338
rect 567234 604338 567266 604894
rect 567822 604338 567854 604894
rect 567234 568894 567854 604338
rect 567234 568338 567266 568894
rect 567822 568338 567854 568894
rect 567234 532894 567854 568338
rect 567234 532338 567266 532894
rect 567822 532338 567854 532894
rect 567234 496894 567854 532338
rect 567234 496338 567266 496894
rect 567822 496338 567854 496894
rect 567234 460894 567854 496338
rect 567234 460338 567266 460894
rect 567822 460338 567854 460894
rect 567234 424894 567854 460338
rect 567234 424338 567266 424894
rect 567822 424338 567854 424894
rect 567234 388894 567854 424338
rect 567234 388338 567266 388894
rect 567822 388338 567854 388894
rect 567234 352894 567854 388338
rect 567234 352338 567266 352894
rect 567822 352338 567854 352894
rect 567234 316894 567854 352338
rect 567234 316338 567266 316894
rect 567822 316338 567854 316894
rect 567234 280894 567854 316338
rect 567234 280338 567266 280894
rect 567822 280338 567854 280894
rect 567234 244894 567854 280338
rect 567234 244338 567266 244894
rect 567822 244338 567854 244894
rect 567234 208894 567854 244338
rect 567234 208338 567266 208894
rect 567822 208338 567854 208894
rect 567234 172894 567854 208338
rect 567234 172338 567266 172894
rect 567822 172338 567854 172894
rect 567234 136894 567854 172338
rect 567234 136338 567266 136894
rect 567822 136338 567854 136894
rect 567234 100894 567854 136338
rect 567234 100338 567266 100894
rect 567822 100338 567854 100894
rect 567234 64894 567854 100338
rect 567234 64338 567266 64894
rect 567822 64338 567854 64894
rect 567234 28894 567854 64338
rect 567234 28338 567266 28894
rect 567822 28338 567854 28894
rect 567234 -5146 567854 28338
rect 567234 -5702 567266 -5146
rect 567822 -5702 567854 -5146
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711002 592062 711558
rect 592618 711002 592650 711558
rect 591070 710598 591690 710630
rect 591070 710042 591102 710598
rect 591658 710042 591690 710598
rect 590110 709638 590730 709670
rect 590110 709082 590142 709638
rect 590698 709082 590730 709638
rect 589150 708678 589770 708710
rect 589150 708122 589182 708678
rect 589738 708122 589770 708678
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707162 588222 707718
rect 588778 707162 588810 707718
rect 581514 706202 581546 706758
rect 582102 706202 582134 706758
rect 570954 680058 570986 680614
rect 571542 680058 571574 680614
rect 570954 644614 571574 680058
rect 570954 644058 570986 644614
rect 571542 644058 571574 644614
rect 570954 608614 571574 644058
rect 570954 608058 570986 608614
rect 571542 608058 571574 608614
rect 570954 572614 571574 608058
rect 570954 572058 570986 572614
rect 571542 572058 571574 572614
rect 570954 536614 571574 572058
rect 570954 536058 570986 536614
rect 571542 536058 571574 536614
rect 570954 500614 571574 536058
rect 570954 500058 570986 500614
rect 571542 500058 571574 500614
rect 570954 464614 571574 500058
rect 570954 464058 570986 464614
rect 571542 464058 571574 464614
rect 570954 428614 571574 464058
rect 570954 428058 570986 428614
rect 571542 428058 571574 428614
rect 570954 392614 571574 428058
rect 570954 392058 570986 392614
rect 571542 392058 571574 392614
rect 570954 356614 571574 392058
rect 570954 356058 570986 356614
rect 571542 356058 571574 356614
rect 570954 320614 571574 356058
rect 570954 320058 570986 320614
rect 571542 320058 571574 320614
rect 570954 284614 571574 320058
rect 570954 284058 570986 284614
rect 571542 284058 571574 284614
rect 570954 248614 571574 284058
rect 570954 248058 570986 248614
rect 571542 248058 571574 248614
rect 570954 212614 571574 248058
rect 570954 212058 570986 212614
rect 571542 212058 571574 212614
rect 570954 176614 571574 212058
rect 570954 176058 570986 176614
rect 571542 176058 571574 176614
rect 570954 140614 571574 176058
rect 570954 140058 570986 140614
rect 571542 140058 571574 140614
rect 570954 104614 571574 140058
rect 570954 104058 570986 104614
rect 571542 104058 571574 104614
rect 570954 68614 571574 104058
rect 570954 68058 570986 68614
rect 571542 68058 571574 68614
rect 570954 32614 571574 68058
rect 570954 32058 570986 32614
rect 571542 32058 571574 32614
rect 552954 -6662 552986 -6106
rect 553542 -6662 553574 -6106
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704282 577826 704838
rect 578382 704282 578414 704838
rect 577794 687454 578414 704282
rect 577794 686898 577826 687454
rect 578382 686898 578414 687454
rect 577794 651454 578414 686898
rect 577794 650898 577826 651454
rect 578382 650898 578414 651454
rect 577794 615454 578414 650898
rect 577794 614898 577826 615454
rect 578382 614898 578414 615454
rect 577794 579454 578414 614898
rect 577794 578898 577826 579454
rect 578382 578898 578414 579454
rect 577794 543454 578414 578898
rect 577794 542898 577826 543454
rect 578382 542898 578414 543454
rect 577794 507454 578414 542898
rect 577794 506898 577826 507454
rect 578382 506898 578414 507454
rect 577794 471454 578414 506898
rect 577794 470898 577826 471454
rect 578382 470898 578414 471454
rect 577794 435454 578414 470898
rect 577794 434898 577826 435454
rect 578382 434898 578414 435454
rect 577794 399454 578414 434898
rect 577794 398898 577826 399454
rect 578382 398898 578414 399454
rect 577794 363454 578414 398898
rect 577794 362898 577826 363454
rect 578382 362898 578414 363454
rect 577794 327454 578414 362898
rect 577794 326898 577826 327454
rect 578382 326898 578414 327454
rect 577794 291454 578414 326898
rect 577794 290898 577826 291454
rect 578382 290898 578414 291454
rect 577794 255454 578414 290898
rect 577794 254898 577826 255454
rect 578382 254898 578414 255454
rect 577794 219454 578414 254898
rect 577794 218898 577826 219454
rect 578382 218898 578414 219454
rect 577794 183454 578414 218898
rect 577794 182898 577826 183454
rect 578382 182898 578414 183454
rect 577794 147454 578414 182898
rect 577794 146898 577826 147454
rect 578382 146898 578414 147454
rect 577794 111454 578414 146898
rect 577794 110898 577826 111454
rect 578382 110898 578414 111454
rect 577794 75454 578414 110898
rect 577794 74898 577826 75454
rect 578382 74898 578414 75454
rect 577794 39454 578414 74898
rect 577794 38898 577826 39454
rect 578382 38898 578414 39454
rect 577794 3454 578414 38898
rect 577794 2898 577826 3454
rect 578382 2898 578414 3454
rect 577794 -346 578414 2898
rect 577794 -902 577826 -346
rect 578382 -902 578414 -346
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706202 587262 706758
rect 587818 706202 587850 706758
rect 586270 705798 586890 705830
rect 586270 705242 586302 705798
rect 586858 705242 586890 705798
rect 581514 690618 581546 691174
rect 582102 690618 582134 691174
rect 581514 655174 582134 690618
rect 581514 654618 581546 655174
rect 582102 654618 582134 655174
rect 581514 619174 582134 654618
rect 581514 618618 581546 619174
rect 582102 618618 582134 619174
rect 581514 583174 582134 618618
rect 581514 582618 581546 583174
rect 582102 582618 582134 583174
rect 581514 547174 582134 582618
rect 581514 546618 581546 547174
rect 582102 546618 582134 547174
rect 581514 511174 582134 546618
rect 581514 510618 581546 511174
rect 582102 510618 582134 511174
rect 581514 475174 582134 510618
rect 581514 474618 581546 475174
rect 582102 474618 582134 475174
rect 581514 439174 582134 474618
rect 581514 438618 581546 439174
rect 582102 438618 582134 439174
rect 581514 403174 582134 438618
rect 581514 402618 581546 403174
rect 582102 402618 582134 403174
rect 581514 367174 582134 402618
rect 581514 366618 581546 367174
rect 582102 366618 582134 367174
rect 581514 331174 582134 366618
rect 581514 330618 581546 331174
rect 582102 330618 582134 331174
rect 581514 295174 582134 330618
rect 581514 294618 581546 295174
rect 582102 294618 582134 295174
rect 581514 259174 582134 294618
rect 581514 258618 581546 259174
rect 582102 258618 582134 259174
rect 581514 223174 582134 258618
rect 581514 222618 581546 223174
rect 582102 222618 582134 223174
rect 581514 187174 582134 222618
rect 581514 186618 581546 187174
rect 582102 186618 582134 187174
rect 581514 151174 582134 186618
rect 581514 150618 581546 151174
rect 582102 150618 582134 151174
rect 581514 115174 582134 150618
rect 581514 114618 581546 115174
rect 582102 114618 582134 115174
rect 581514 79174 582134 114618
rect 581514 78618 581546 79174
rect 582102 78618 582134 79174
rect 581514 43174 582134 78618
rect 581514 42618 581546 43174
rect 582102 42618 582134 43174
rect 581514 7174 582134 42618
rect 581514 6618 581546 7174
rect 582102 6618 582134 7174
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704282 585342 704838
rect 585898 704282 585930 704838
rect 585310 687454 585930 704282
rect 585310 686898 585342 687454
rect 585898 686898 585930 687454
rect 585310 651454 585930 686898
rect 585310 650898 585342 651454
rect 585898 650898 585930 651454
rect 585310 615454 585930 650898
rect 585310 614898 585342 615454
rect 585898 614898 585930 615454
rect 585310 579454 585930 614898
rect 585310 578898 585342 579454
rect 585898 578898 585930 579454
rect 585310 543454 585930 578898
rect 585310 542898 585342 543454
rect 585898 542898 585930 543454
rect 585310 507454 585930 542898
rect 585310 506898 585342 507454
rect 585898 506898 585930 507454
rect 585310 471454 585930 506898
rect 585310 470898 585342 471454
rect 585898 470898 585930 471454
rect 585310 435454 585930 470898
rect 585310 434898 585342 435454
rect 585898 434898 585930 435454
rect 585310 399454 585930 434898
rect 585310 398898 585342 399454
rect 585898 398898 585930 399454
rect 585310 363454 585930 398898
rect 585310 362898 585342 363454
rect 585898 362898 585930 363454
rect 585310 327454 585930 362898
rect 585310 326898 585342 327454
rect 585898 326898 585930 327454
rect 585310 291454 585930 326898
rect 585310 290898 585342 291454
rect 585898 290898 585930 291454
rect 585310 255454 585930 290898
rect 585310 254898 585342 255454
rect 585898 254898 585930 255454
rect 585310 219454 585930 254898
rect 585310 218898 585342 219454
rect 585898 218898 585930 219454
rect 585310 183454 585930 218898
rect 585310 182898 585342 183454
rect 585898 182898 585930 183454
rect 585310 147454 585930 182898
rect 585310 146898 585342 147454
rect 585898 146898 585930 147454
rect 585310 111454 585930 146898
rect 585310 110898 585342 111454
rect 585898 110898 585930 111454
rect 585310 75454 585930 110898
rect 585310 74898 585342 75454
rect 585898 74898 585930 75454
rect 585310 39454 585930 74898
rect 585310 38898 585342 39454
rect 585898 38898 585930 39454
rect 585310 3454 585930 38898
rect 585310 2898 585342 3454
rect 585898 2898 585930 3454
rect 585310 -346 585930 2898
rect 585310 -902 585342 -346
rect 585898 -902 585930 -346
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 668898 586302 669454
rect 586858 668898 586890 669454
rect 586270 633454 586890 668898
rect 586270 632898 586302 633454
rect 586858 632898 586890 633454
rect 586270 597454 586890 632898
rect 586270 596898 586302 597454
rect 586858 596898 586890 597454
rect 586270 561454 586890 596898
rect 586270 560898 586302 561454
rect 586858 560898 586890 561454
rect 586270 525454 586890 560898
rect 586270 524898 586302 525454
rect 586858 524898 586890 525454
rect 586270 489454 586890 524898
rect 586270 488898 586302 489454
rect 586858 488898 586890 489454
rect 586270 453454 586890 488898
rect 586270 452898 586302 453454
rect 586858 452898 586890 453454
rect 586270 417454 586890 452898
rect 586270 416898 586302 417454
rect 586858 416898 586890 417454
rect 586270 381454 586890 416898
rect 586270 380898 586302 381454
rect 586858 380898 586890 381454
rect 586270 345454 586890 380898
rect 586270 344898 586302 345454
rect 586858 344898 586890 345454
rect 586270 309454 586890 344898
rect 586270 308898 586302 309454
rect 586858 308898 586890 309454
rect 586270 273454 586890 308898
rect 586270 272898 586302 273454
rect 586858 272898 586890 273454
rect 586270 237454 586890 272898
rect 586270 236898 586302 237454
rect 586858 236898 586890 237454
rect 586270 201454 586890 236898
rect 586270 200898 586302 201454
rect 586858 200898 586890 201454
rect 586270 165454 586890 200898
rect 586270 164898 586302 165454
rect 586858 164898 586890 165454
rect 586270 129454 586890 164898
rect 586270 128898 586302 129454
rect 586858 128898 586890 129454
rect 586270 93454 586890 128898
rect 586270 92898 586302 93454
rect 586858 92898 586890 93454
rect 586270 57454 586890 92898
rect 586270 56898 586302 57454
rect 586858 56898 586890 57454
rect 586270 21454 586890 56898
rect 586270 20898 586302 21454
rect 586858 20898 586890 21454
rect 586270 -1306 586890 20898
rect 586270 -1862 586302 -1306
rect 586858 -1862 586890 -1306
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690618 587262 691174
rect 587818 690618 587850 691174
rect 587230 655174 587850 690618
rect 587230 654618 587262 655174
rect 587818 654618 587850 655174
rect 587230 619174 587850 654618
rect 587230 618618 587262 619174
rect 587818 618618 587850 619174
rect 587230 583174 587850 618618
rect 587230 582618 587262 583174
rect 587818 582618 587850 583174
rect 587230 547174 587850 582618
rect 587230 546618 587262 547174
rect 587818 546618 587850 547174
rect 587230 511174 587850 546618
rect 587230 510618 587262 511174
rect 587818 510618 587850 511174
rect 587230 475174 587850 510618
rect 587230 474618 587262 475174
rect 587818 474618 587850 475174
rect 587230 439174 587850 474618
rect 587230 438618 587262 439174
rect 587818 438618 587850 439174
rect 587230 403174 587850 438618
rect 587230 402618 587262 403174
rect 587818 402618 587850 403174
rect 587230 367174 587850 402618
rect 587230 366618 587262 367174
rect 587818 366618 587850 367174
rect 587230 331174 587850 366618
rect 587230 330618 587262 331174
rect 587818 330618 587850 331174
rect 587230 295174 587850 330618
rect 587230 294618 587262 295174
rect 587818 294618 587850 295174
rect 587230 259174 587850 294618
rect 587230 258618 587262 259174
rect 587818 258618 587850 259174
rect 587230 223174 587850 258618
rect 587230 222618 587262 223174
rect 587818 222618 587850 223174
rect 587230 187174 587850 222618
rect 587230 186618 587262 187174
rect 587818 186618 587850 187174
rect 587230 151174 587850 186618
rect 587230 150618 587262 151174
rect 587818 150618 587850 151174
rect 587230 115174 587850 150618
rect 587230 114618 587262 115174
rect 587818 114618 587850 115174
rect 587230 79174 587850 114618
rect 587230 78618 587262 79174
rect 587818 78618 587850 79174
rect 587230 43174 587850 78618
rect 587230 42618 587262 43174
rect 587818 42618 587850 43174
rect 587230 7174 587850 42618
rect 587230 6618 587262 7174
rect 587818 6618 587850 7174
rect 581514 -2822 581546 -2266
rect 582102 -2822 582134 -2266
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2822 587262 -2266
rect 587818 -2822 587850 -2266
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672618 588222 673174
rect 588778 672618 588810 673174
rect 588190 637174 588810 672618
rect 588190 636618 588222 637174
rect 588778 636618 588810 637174
rect 588190 601174 588810 636618
rect 588190 600618 588222 601174
rect 588778 600618 588810 601174
rect 588190 565174 588810 600618
rect 588190 564618 588222 565174
rect 588778 564618 588810 565174
rect 588190 529174 588810 564618
rect 588190 528618 588222 529174
rect 588778 528618 588810 529174
rect 588190 493174 588810 528618
rect 588190 492618 588222 493174
rect 588778 492618 588810 493174
rect 588190 457174 588810 492618
rect 588190 456618 588222 457174
rect 588778 456618 588810 457174
rect 588190 421174 588810 456618
rect 588190 420618 588222 421174
rect 588778 420618 588810 421174
rect 588190 385174 588810 420618
rect 588190 384618 588222 385174
rect 588778 384618 588810 385174
rect 588190 349174 588810 384618
rect 588190 348618 588222 349174
rect 588778 348618 588810 349174
rect 588190 313174 588810 348618
rect 588190 312618 588222 313174
rect 588778 312618 588810 313174
rect 588190 277174 588810 312618
rect 588190 276618 588222 277174
rect 588778 276618 588810 277174
rect 588190 241174 588810 276618
rect 588190 240618 588222 241174
rect 588778 240618 588810 241174
rect 588190 205174 588810 240618
rect 588190 204618 588222 205174
rect 588778 204618 588810 205174
rect 588190 169174 588810 204618
rect 588190 168618 588222 169174
rect 588778 168618 588810 169174
rect 588190 133174 588810 168618
rect 588190 132618 588222 133174
rect 588778 132618 588810 133174
rect 588190 97174 588810 132618
rect 588190 96618 588222 97174
rect 588778 96618 588810 97174
rect 588190 61174 588810 96618
rect 588190 60618 588222 61174
rect 588778 60618 588810 61174
rect 588190 25174 588810 60618
rect 588190 24618 588222 25174
rect 588778 24618 588810 25174
rect 588190 -3226 588810 24618
rect 588190 -3782 588222 -3226
rect 588778 -3782 588810 -3226
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694338 589182 694894
rect 589738 694338 589770 694894
rect 589150 658894 589770 694338
rect 589150 658338 589182 658894
rect 589738 658338 589770 658894
rect 589150 622894 589770 658338
rect 589150 622338 589182 622894
rect 589738 622338 589770 622894
rect 589150 586894 589770 622338
rect 589150 586338 589182 586894
rect 589738 586338 589770 586894
rect 589150 550894 589770 586338
rect 589150 550338 589182 550894
rect 589738 550338 589770 550894
rect 589150 514894 589770 550338
rect 589150 514338 589182 514894
rect 589738 514338 589770 514894
rect 589150 478894 589770 514338
rect 589150 478338 589182 478894
rect 589738 478338 589770 478894
rect 589150 442894 589770 478338
rect 589150 442338 589182 442894
rect 589738 442338 589770 442894
rect 589150 406894 589770 442338
rect 589150 406338 589182 406894
rect 589738 406338 589770 406894
rect 589150 370894 589770 406338
rect 589150 370338 589182 370894
rect 589738 370338 589770 370894
rect 589150 334894 589770 370338
rect 589150 334338 589182 334894
rect 589738 334338 589770 334894
rect 589150 298894 589770 334338
rect 589150 298338 589182 298894
rect 589738 298338 589770 298894
rect 589150 262894 589770 298338
rect 589150 262338 589182 262894
rect 589738 262338 589770 262894
rect 589150 226894 589770 262338
rect 589150 226338 589182 226894
rect 589738 226338 589770 226894
rect 589150 190894 589770 226338
rect 589150 190338 589182 190894
rect 589738 190338 589770 190894
rect 589150 154894 589770 190338
rect 589150 154338 589182 154894
rect 589738 154338 589770 154894
rect 589150 118894 589770 154338
rect 589150 118338 589182 118894
rect 589738 118338 589770 118894
rect 589150 82894 589770 118338
rect 589150 82338 589182 82894
rect 589738 82338 589770 82894
rect 589150 46894 589770 82338
rect 589150 46338 589182 46894
rect 589738 46338 589770 46894
rect 589150 10894 589770 46338
rect 589150 10338 589182 10894
rect 589738 10338 589770 10894
rect 589150 -4186 589770 10338
rect 589150 -4742 589182 -4186
rect 589738 -4742 589770 -4186
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676338 590142 676894
rect 590698 676338 590730 676894
rect 590110 640894 590730 676338
rect 590110 640338 590142 640894
rect 590698 640338 590730 640894
rect 590110 604894 590730 640338
rect 590110 604338 590142 604894
rect 590698 604338 590730 604894
rect 590110 568894 590730 604338
rect 590110 568338 590142 568894
rect 590698 568338 590730 568894
rect 590110 532894 590730 568338
rect 590110 532338 590142 532894
rect 590698 532338 590730 532894
rect 590110 496894 590730 532338
rect 590110 496338 590142 496894
rect 590698 496338 590730 496894
rect 590110 460894 590730 496338
rect 590110 460338 590142 460894
rect 590698 460338 590730 460894
rect 590110 424894 590730 460338
rect 590110 424338 590142 424894
rect 590698 424338 590730 424894
rect 590110 388894 590730 424338
rect 590110 388338 590142 388894
rect 590698 388338 590730 388894
rect 590110 352894 590730 388338
rect 590110 352338 590142 352894
rect 590698 352338 590730 352894
rect 590110 316894 590730 352338
rect 590110 316338 590142 316894
rect 590698 316338 590730 316894
rect 590110 280894 590730 316338
rect 590110 280338 590142 280894
rect 590698 280338 590730 280894
rect 590110 244894 590730 280338
rect 590110 244338 590142 244894
rect 590698 244338 590730 244894
rect 590110 208894 590730 244338
rect 590110 208338 590142 208894
rect 590698 208338 590730 208894
rect 590110 172894 590730 208338
rect 590110 172338 590142 172894
rect 590698 172338 590730 172894
rect 590110 136894 590730 172338
rect 590110 136338 590142 136894
rect 590698 136338 590730 136894
rect 590110 100894 590730 136338
rect 590110 100338 590142 100894
rect 590698 100338 590730 100894
rect 590110 64894 590730 100338
rect 590110 64338 590142 64894
rect 590698 64338 590730 64894
rect 590110 28894 590730 64338
rect 590110 28338 590142 28894
rect 590698 28338 590730 28894
rect 590110 -5146 590730 28338
rect 590110 -5702 590142 -5146
rect 590698 -5702 590730 -5146
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698058 591102 698614
rect 591658 698058 591690 698614
rect 591070 662614 591690 698058
rect 591070 662058 591102 662614
rect 591658 662058 591690 662614
rect 591070 626614 591690 662058
rect 591070 626058 591102 626614
rect 591658 626058 591690 626614
rect 591070 590614 591690 626058
rect 591070 590058 591102 590614
rect 591658 590058 591690 590614
rect 591070 554614 591690 590058
rect 591070 554058 591102 554614
rect 591658 554058 591690 554614
rect 591070 518614 591690 554058
rect 591070 518058 591102 518614
rect 591658 518058 591690 518614
rect 591070 482614 591690 518058
rect 591070 482058 591102 482614
rect 591658 482058 591690 482614
rect 591070 446614 591690 482058
rect 591070 446058 591102 446614
rect 591658 446058 591690 446614
rect 591070 410614 591690 446058
rect 591070 410058 591102 410614
rect 591658 410058 591690 410614
rect 591070 374614 591690 410058
rect 591070 374058 591102 374614
rect 591658 374058 591690 374614
rect 591070 338614 591690 374058
rect 591070 338058 591102 338614
rect 591658 338058 591690 338614
rect 591070 302614 591690 338058
rect 591070 302058 591102 302614
rect 591658 302058 591690 302614
rect 591070 266614 591690 302058
rect 591070 266058 591102 266614
rect 591658 266058 591690 266614
rect 591070 230614 591690 266058
rect 591070 230058 591102 230614
rect 591658 230058 591690 230614
rect 591070 194614 591690 230058
rect 591070 194058 591102 194614
rect 591658 194058 591690 194614
rect 591070 158614 591690 194058
rect 591070 158058 591102 158614
rect 591658 158058 591690 158614
rect 591070 122614 591690 158058
rect 591070 122058 591102 122614
rect 591658 122058 591690 122614
rect 591070 86614 591690 122058
rect 591070 86058 591102 86614
rect 591658 86058 591690 86614
rect 591070 50614 591690 86058
rect 591070 50058 591102 50614
rect 591658 50058 591690 50614
rect 591070 14614 591690 50058
rect 591070 14058 591102 14614
rect 591658 14058 591690 14614
rect 591070 -6106 591690 14058
rect 591070 -6662 591102 -6106
rect 591658 -6662 591690 -6106
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680058 592062 680614
rect 592618 680058 592650 680614
rect 592030 644614 592650 680058
rect 592030 644058 592062 644614
rect 592618 644058 592650 644614
rect 592030 608614 592650 644058
rect 592030 608058 592062 608614
rect 592618 608058 592650 608614
rect 592030 572614 592650 608058
rect 592030 572058 592062 572614
rect 592618 572058 592650 572614
rect 592030 536614 592650 572058
rect 592030 536058 592062 536614
rect 592618 536058 592650 536614
rect 592030 500614 592650 536058
rect 592030 500058 592062 500614
rect 592618 500058 592650 500614
rect 592030 464614 592650 500058
rect 592030 464058 592062 464614
rect 592618 464058 592650 464614
rect 592030 428614 592650 464058
rect 592030 428058 592062 428614
rect 592618 428058 592650 428614
rect 592030 392614 592650 428058
rect 592030 392058 592062 392614
rect 592618 392058 592650 392614
rect 592030 356614 592650 392058
rect 592030 356058 592062 356614
rect 592618 356058 592650 356614
rect 592030 320614 592650 356058
rect 592030 320058 592062 320614
rect 592618 320058 592650 320614
rect 592030 284614 592650 320058
rect 592030 284058 592062 284614
rect 592618 284058 592650 284614
rect 592030 248614 592650 284058
rect 592030 248058 592062 248614
rect 592618 248058 592650 248614
rect 592030 212614 592650 248058
rect 592030 212058 592062 212614
rect 592618 212058 592650 212614
rect 592030 176614 592650 212058
rect 592030 176058 592062 176614
rect 592618 176058 592650 176614
rect 592030 140614 592650 176058
rect 592030 140058 592062 140614
rect 592618 140058 592650 140614
rect 592030 104614 592650 140058
rect 592030 104058 592062 104614
rect 592618 104058 592650 104614
rect 592030 68614 592650 104058
rect 592030 68058 592062 68614
rect 592618 68058 592650 68614
rect 592030 32614 592650 68058
rect 592030 32058 592062 32614
rect 592618 32058 592650 32614
rect 570954 -7622 570986 -7066
rect 571542 -7622 571574 -7066
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7622 592062 -7066
rect 592618 -7622 592650 -7066
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711002 -8138 711558
rect -8694 680058 -8138 680614
rect -8694 644058 -8138 644614
rect -8694 608058 -8138 608614
rect -8694 572058 -8138 572614
rect -8694 536058 -8138 536614
rect -8694 500058 -8138 500614
rect -8694 464058 -8138 464614
rect -8694 428058 -8138 428614
rect -8694 392058 -8138 392614
rect -8694 356058 -8138 356614
rect -8694 320058 -8138 320614
rect -8694 284058 -8138 284614
rect -8694 248058 -8138 248614
rect -8694 212058 -8138 212614
rect -8694 176058 -8138 176614
rect -8694 140058 -8138 140614
rect -8694 104058 -8138 104614
rect -8694 68058 -8138 68614
rect -8694 32058 -8138 32614
rect -7734 710042 -7178 710598
rect 12986 710042 13542 710598
rect -7734 698058 -7178 698614
rect -7734 662058 -7178 662614
rect -7734 626058 -7178 626614
rect -7734 590058 -7178 590614
rect -7734 554058 -7178 554614
rect -7734 518058 -7178 518614
rect -7734 482058 -7178 482614
rect -7734 446058 -7178 446614
rect -7734 410058 -7178 410614
rect -7734 374058 -7178 374614
rect -7734 338058 -7178 338614
rect -7734 302058 -7178 302614
rect -7734 266058 -7178 266614
rect -7734 230058 -7178 230614
rect -7734 194058 -7178 194614
rect -7734 158058 -7178 158614
rect -7734 122058 -7178 122614
rect -7734 86058 -7178 86614
rect -7734 50058 -7178 50614
rect -7734 14058 -7178 14614
rect -6774 709082 -6218 709638
rect -6774 676338 -6218 676894
rect -6774 640338 -6218 640894
rect -6774 604338 -6218 604894
rect -6774 568338 -6218 568894
rect -6774 532338 -6218 532894
rect -6774 496338 -6218 496894
rect -6774 460338 -6218 460894
rect -6774 424338 -6218 424894
rect -6774 388338 -6218 388894
rect -6774 352338 -6218 352894
rect -6774 316338 -6218 316894
rect -6774 280338 -6218 280894
rect -6774 244338 -6218 244894
rect -6774 208338 -6218 208894
rect -6774 172338 -6218 172894
rect -6774 136338 -6218 136894
rect -6774 100338 -6218 100894
rect -6774 64338 -6218 64894
rect -6774 28338 -6218 28894
rect -5814 708122 -5258 708678
rect 9266 708122 9822 708678
rect -5814 694338 -5258 694894
rect -5814 658338 -5258 658894
rect -5814 622338 -5258 622894
rect -5814 586338 -5258 586894
rect -5814 550338 -5258 550894
rect -5814 514338 -5258 514894
rect -5814 478338 -5258 478894
rect -5814 442338 -5258 442894
rect -5814 406338 -5258 406894
rect -5814 370338 -5258 370894
rect -5814 334338 -5258 334894
rect -5814 298338 -5258 298894
rect -5814 262338 -5258 262894
rect -5814 226338 -5258 226894
rect -5814 190338 -5258 190894
rect -5814 154338 -5258 154894
rect -5814 118338 -5258 118894
rect -5814 82338 -5258 82894
rect -5814 46338 -5258 46894
rect -5814 10338 -5258 10894
rect -4854 707162 -4298 707718
rect -4854 672618 -4298 673174
rect -4854 636618 -4298 637174
rect -4854 600618 -4298 601174
rect -4854 564618 -4298 565174
rect -4854 528618 -4298 529174
rect -4854 492618 -4298 493174
rect -4854 456618 -4298 457174
rect -4854 420618 -4298 421174
rect -4854 384618 -4298 385174
rect -4854 348618 -4298 349174
rect -4854 312618 -4298 313174
rect -4854 276618 -4298 277174
rect -4854 240618 -4298 241174
rect -4854 204618 -4298 205174
rect -4854 168618 -4298 169174
rect -4854 132618 -4298 133174
rect -4854 96618 -4298 97174
rect -4854 60618 -4298 61174
rect -4854 24618 -4298 25174
rect -3894 706202 -3338 706758
rect 5546 706202 6102 706758
rect -3894 690618 -3338 691174
rect -3894 654618 -3338 655174
rect -3894 618618 -3338 619174
rect -3894 582618 -3338 583174
rect -3894 546618 -3338 547174
rect -3894 510618 -3338 511174
rect -3894 474618 -3338 475174
rect -3894 438618 -3338 439174
rect -3894 402618 -3338 403174
rect -3894 366618 -3338 367174
rect -3894 330618 -3338 331174
rect -3894 294618 -3338 295174
rect -3894 258618 -3338 259174
rect -3894 222618 -3338 223174
rect -3894 186618 -3338 187174
rect -3894 150618 -3338 151174
rect -3894 114618 -3338 115174
rect -3894 78618 -3338 79174
rect -3894 42618 -3338 43174
rect -3894 6618 -3338 7174
rect -2934 705242 -2378 705798
rect -2934 668898 -2378 669454
rect -2934 632898 -2378 633454
rect -2934 596898 -2378 597454
rect -2934 560898 -2378 561454
rect -2934 524898 -2378 525454
rect -2934 488898 -2378 489454
rect -2934 452898 -2378 453454
rect -2934 416898 -2378 417454
rect -2934 380898 -2378 381454
rect -2934 344898 -2378 345454
rect -2934 308898 -2378 309454
rect -2934 272898 -2378 273454
rect -2934 236898 -2378 237454
rect -2934 200898 -2378 201454
rect -2934 164898 -2378 165454
rect -2934 128898 -2378 129454
rect -2934 92898 -2378 93454
rect -2934 56898 -2378 57454
rect -2934 20898 -2378 21454
rect -1974 704282 -1418 704838
rect -1974 686898 -1418 687454
rect -1974 650898 -1418 651454
rect -1974 614898 -1418 615454
rect -1974 578898 -1418 579454
rect -1974 542898 -1418 543454
rect -1974 506898 -1418 507454
rect -1974 470898 -1418 471454
rect -1974 434898 -1418 435454
rect -1974 398898 -1418 399454
rect -1974 362898 -1418 363454
rect -1974 326898 -1418 327454
rect -1974 290898 -1418 291454
rect -1974 254898 -1418 255454
rect -1974 218898 -1418 219454
rect -1974 182898 -1418 183454
rect -1974 146898 -1418 147454
rect -1974 110898 -1418 111454
rect -1974 74898 -1418 75454
rect -1974 38898 -1418 39454
rect -1974 2898 -1418 3454
rect -1974 -902 -1418 -346
rect 1826 704282 2382 704838
rect 1826 686898 2382 687454
rect 1826 650898 2382 651454
rect 1826 614898 2382 615454
rect 1826 578898 2382 579454
rect 1826 542898 2382 543454
rect 1826 506898 2382 507454
rect 1826 470898 2382 471454
rect 1826 434898 2382 435454
rect 1826 398898 2382 399454
rect 1826 362898 2382 363454
rect 1826 326898 2382 327454
rect 1826 290898 2382 291454
rect 1826 254898 2382 255454
rect 1826 218898 2382 219454
rect 1826 182898 2382 183454
rect 1826 146898 2382 147454
rect 1826 110898 2382 111454
rect 1826 74898 2382 75454
rect 1826 38898 2382 39454
rect 1826 2898 2382 3454
rect 1826 -902 2382 -346
rect -2934 -1862 -2378 -1306
rect 5546 690618 6102 691174
rect 5546 654618 6102 655174
rect 5546 618618 6102 619174
rect 5546 582618 6102 583174
rect 5546 546618 6102 547174
rect 5546 510618 6102 511174
rect 5546 474618 6102 475174
rect 5546 438618 6102 439174
rect 5546 402618 6102 403174
rect 5546 366618 6102 367174
rect 5546 330618 6102 331174
rect 5546 294618 6102 295174
rect 5546 258618 6102 259174
rect 5546 222618 6102 223174
rect 5546 186618 6102 187174
rect 5546 150618 6102 151174
rect 5546 114618 6102 115174
rect 5546 78618 6102 79174
rect 5546 42618 6102 43174
rect 5546 6618 6102 7174
rect -3894 -2822 -3338 -2266
rect 5546 -2822 6102 -2266
rect -4854 -3782 -4298 -3226
rect 9266 694338 9822 694894
rect 9266 658338 9822 658894
rect 9266 622338 9822 622894
rect 9266 586338 9822 586894
rect 9266 550338 9822 550894
rect 9266 514338 9822 514894
rect 9266 478338 9822 478894
rect 9266 442338 9822 442894
rect 9266 406338 9822 406894
rect 9266 370338 9822 370894
rect 9266 334338 9822 334894
rect 9266 298338 9822 298894
rect 9266 262338 9822 262894
rect 9266 226338 9822 226894
rect 9266 190338 9822 190894
rect 9266 154338 9822 154894
rect 9266 118338 9822 118894
rect 9266 82338 9822 82894
rect 9266 46338 9822 46894
rect 9266 10338 9822 10894
rect -5814 -4742 -5258 -4186
rect 9266 -4742 9822 -4186
rect -6774 -5702 -6218 -5146
rect 30986 711002 31542 711558
rect 27266 709082 27822 709638
rect 23546 707162 24102 707718
rect 12986 698058 13542 698614
rect 12986 662058 13542 662614
rect 12986 626058 13542 626614
rect 12986 590058 13542 590614
rect 12986 554058 13542 554614
rect 12986 518058 13542 518614
rect 12986 482058 13542 482614
rect 12986 446058 13542 446614
rect 12986 410058 13542 410614
rect 12986 374058 13542 374614
rect 12986 338058 13542 338614
rect 12986 302058 13542 302614
rect 12986 266058 13542 266614
rect 12986 230058 13542 230614
rect 12986 194058 13542 194614
rect 12986 158058 13542 158614
rect 12986 122058 13542 122614
rect 12986 86058 13542 86614
rect 12986 50058 13542 50614
rect 12986 14058 13542 14614
rect -7734 -6662 -7178 -6106
rect 19826 705242 20382 705798
rect 19826 668898 20382 669454
rect 19826 632898 20382 633454
rect 19826 596898 20382 597454
rect 19826 560898 20382 561454
rect 19826 524898 20382 525454
rect 19826 488898 20382 489454
rect 19826 452898 20382 453454
rect 19826 416898 20382 417454
rect 19826 380898 20382 381454
rect 19826 344898 20382 345454
rect 19826 308898 20382 309454
rect 19826 272898 20382 273454
rect 19826 236898 20382 237454
rect 19826 200898 20382 201454
rect 19826 164898 20382 165454
rect 19826 128898 20382 129454
rect 19826 92898 20382 93454
rect 19826 56898 20382 57454
rect 19826 20898 20382 21454
rect 19826 -1862 20382 -1306
rect 23546 672618 24102 673174
rect 23546 636618 24102 637174
rect 23546 600618 24102 601174
rect 23546 564618 24102 565174
rect 23546 528618 24102 529174
rect 23546 492618 24102 493174
rect 23546 456618 24102 457174
rect 23546 420618 24102 421174
rect 23546 384618 24102 385174
rect 23546 348618 24102 349174
rect 23546 312618 24102 313174
rect 23546 276618 24102 277174
rect 23546 240618 24102 241174
rect 23546 204618 24102 205174
rect 23546 168618 24102 169174
rect 23546 132618 24102 133174
rect 23546 96618 24102 97174
rect 23546 60618 24102 61174
rect 23546 24618 24102 25174
rect 23546 -3782 24102 -3226
rect 27266 676338 27822 676894
rect 27266 640338 27822 640894
rect 27266 604338 27822 604894
rect 27266 568338 27822 568894
rect 27266 532338 27822 532894
rect 27266 496338 27822 496894
rect 27266 460338 27822 460894
rect 27266 424338 27822 424894
rect 27266 388338 27822 388894
rect 27266 352338 27822 352894
rect 27266 316338 27822 316894
rect 27266 280338 27822 280894
rect 27266 244338 27822 244894
rect 27266 208338 27822 208894
rect 27266 172338 27822 172894
rect 27266 136338 27822 136894
rect 27266 100338 27822 100894
rect 27266 64338 27822 64894
rect 27266 28338 27822 28894
rect 27266 -5702 27822 -5146
rect 48986 710042 49542 710598
rect 45266 708122 45822 708678
rect 41546 706202 42102 706758
rect 30986 680058 31542 680614
rect 30986 644058 31542 644614
rect 30986 608058 31542 608614
rect 30986 572058 31542 572614
rect 30986 536058 31542 536614
rect 30986 500058 31542 500614
rect 30986 464058 31542 464614
rect 30986 428058 31542 428614
rect 30986 392058 31542 392614
rect 30986 356058 31542 356614
rect 30986 320058 31542 320614
rect 30986 284058 31542 284614
rect 30986 248058 31542 248614
rect 30986 212058 31542 212614
rect 30986 176058 31542 176614
rect 30986 140058 31542 140614
rect 30986 104058 31542 104614
rect 30986 68058 31542 68614
rect 30986 32058 31542 32614
rect 12986 -6662 13542 -6106
rect -8694 -7622 -8138 -7066
rect 37826 704282 38382 704838
rect 37826 686898 38382 687454
rect 37826 650898 38382 651454
rect 37826 614898 38382 615454
rect 37826 578898 38382 579454
rect 37826 542898 38382 543454
rect 37826 506898 38382 507454
rect 37826 470898 38382 471454
rect 37826 434898 38382 435454
rect 37826 398898 38382 399454
rect 37826 362898 38382 363454
rect 37826 326898 38382 327454
rect 37826 290898 38382 291454
rect 37826 254898 38382 255454
rect 37826 218898 38382 219454
rect 37826 182898 38382 183454
rect 37826 146898 38382 147454
rect 37826 110898 38382 111454
rect 37826 74898 38382 75454
rect 37826 38898 38382 39454
rect 37826 2898 38382 3454
rect 37826 -902 38382 -346
rect 41546 690618 42102 691174
rect 41546 654618 42102 655174
rect 41546 618618 42102 619174
rect 41546 582618 42102 583174
rect 41546 546618 42102 547174
rect 41546 510618 42102 511174
rect 41546 474618 42102 475174
rect 41546 438618 42102 439174
rect 41546 402618 42102 403174
rect 41546 366618 42102 367174
rect 41546 330618 42102 331174
rect 41546 294618 42102 295174
rect 41546 258618 42102 259174
rect 41546 222618 42102 223174
rect 41546 186618 42102 187174
rect 41546 150618 42102 151174
rect 41546 114618 42102 115174
rect 41546 78618 42102 79174
rect 41546 42618 42102 43174
rect 41546 6618 42102 7174
rect 41546 -2822 42102 -2266
rect 45266 694338 45822 694894
rect 45266 658338 45822 658894
rect 45266 622338 45822 622894
rect 45266 586338 45822 586894
rect 45266 550338 45822 550894
rect 45266 514338 45822 514894
rect 45266 478338 45822 478894
rect 45266 442338 45822 442894
rect 45266 406338 45822 406894
rect 45266 370338 45822 370894
rect 45266 334338 45822 334894
rect 45266 298338 45822 298894
rect 45266 262338 45822 262894
rect 45266 226338 45822 226894
rect 45266 190338 45822 190894
rect 45266 154338 45822 154894
rect 45266 118338 45822 118894
rect 45266 82338 45822 82894
rect 45266 46338 45822 46894
rect 45266 10338 45822 10894
rect 45266 -4742 45822 -4186
rect 66986 711002 67542 711558
rect 63266 709082 63822 709638
rect 59546 707162 60102 707718
rect 48986 698058 49542 698614
rect 48986 662058 49542 662614
rect 48986 626058 49542 626614
rect 48986 590058 49542 590614
rect 48986 554058 49542 554614
rect 48986 518058 49542 518614
rect 48986 482058 49542 482614
rect 48986 446058 49542 446614
rect 48986 410058 49542 410614
rect 48986 374058 49542 374614
rect 48986 338058 49542 338614
rect 48986 302058 49542 302614
rect 48986 266058 49542 266614
rect 48986 230058 49542 230614
rect 48986 194058 49542 194614
rect 48986 158058 49542 158614
rect 48986 122058 49542 122614
rect 48986 86058 49542 86614
rect 48986 50058 49542 50614
rect 48986 14058 49542 14614
rect 30986 -7622 31542 -7066
rect 55826 705242 56382 705798
rect 55826 668898 56382 669454
rect 55826 632898 56382 633454
rect 55826 596898 56382 597454
rect 55826 560898 56382 561454
rect 55826 524898 56382 525454
rect 55826 488898 56382 489454
rect 55826 452898 56382 453454
rect 55826 416898 56382 417454
rect 55826 380898 56382 381454
rect 55826 344898 56382 345454
rect 55826 308898 56382 309454
rect 55826 272898 56382 273454
rect 55826 236898 56382 237454
rect 55826 200898 56382 201454
rect 55826 164898 56382 165454
rect 55826 128898 56382 129454
rect 55826 92898 56382 93454
rect 55826 56898 56382 57454
rect 55826 20898 56382 21454
rect 55826 -1862 56382 -1306
rect 59546 672618 60102 673174
rect 59546 636618 60102 637174
rect 59546 600618 60102 601174
rect 59546 564618 60102 565174
rect 59546 528618 60102 529174
rect 59546 492618 60102 493174
rect 59546 456618 60102 457174
rect 59546 420618 60102 421174
rect 59546 384618 60102 385174
rect 59546 348618 60102 349174
rect 59546 312618 60102 313174
rect 59546 276618 60102 277174
rect 59546 240618 60102 241174
rect 59546 204618 60102 205174
rect 59546 168618 60102 169174
rect 59546 132618 60102 133174
rect 59546 96618 60102 97174
rect 59546 60618 60102 61174
rect 59546 24618 60102 25174
rect 59546 -3782 60102 -3226
rect 63266 676338 63822 676894
rect 63266 640338 63822 640894
rect 63266 604338 63822 604894
rect 63266 568338 63822 568894
rect 63266 532338 63822 532894
rect 63266 496338 63822 496894
rect 63266 460338 63822 460894
rect 63266 424338 63822 424894
rect 63266 388338 63822 388894
rect 63266 352338 63822 352894
rect 63266 316338 63822 316894
rect 63266 280338 63822 280894
rect 63266 244338 63822 244894
rect 63266 208338 63822 208894
rect 63266 172338 63822 172894
rect 63266 136338 63822 136894
rect 63266 100338 63822 100894
rect 63266 64338 63822 64894
rect 63266 28338 63822 28894
rect 63266 -5702 63822 -5146
rect 84986 710042 85542 710598
rect 81266 708122 81822 708678
rect 77546 706202 78102 706758
rect 66986 680058 67542 680614
rect 66986 644058 67542 644614
rect 66986 608058 67542 608614
rect 66986 572058 67542 572614
rect 66986 536058 67542 536614
rect 66986 500058 67542 500614
rect 66986 464058 67542 464614
rect 66986 428058 67542 428614
rect 66986 392058 67542 392614
rect 66986 356058 67542 356614
rect 66986 320058 67542 320614
rect 66986 284058 67542 284614
rect 66986 248058 67542 248614
rect 66986 212058 67542 212614
rect 66986 176058 67542 176614
rect 66986 140058 67542 140614
rect 66986 104058 67542 104614
rect 66986 68058 67542 68614
rect 66986 32058 67542 32614
rect 48986 -6662 49542 -6106
rect 73826 704282 74382 704838
rect 73826 686898 74382 687454
rect 73826 650898 74382 651454
rect 73826 614898 74382 615454
rect 73826 578898 74382 579454
rect 73826 542898 74382 543454
rect 73826 506898 74382 507454
rect 73826 470898 74382 471454
rect 73826 434898 74382 435454
rect 73826 398898 74382 399454
rect 73826 362898 74382 363454
rect 73826 326898 74382 327454
rect 73826 290898 74382 291454
rect 73826 254898 74382 255454
rect 73826 218898 74382 219454
rect 73826 182898 74382 183454
rect 73826 146898 74382 147454
rect 73826 110898 74382 111454
rect 73826 74898 74382 75454
rect 73826 38898 74382 39454
rect 73826 2898 74382 3454
rect 73826 -902 74382 -346
rect 77546 690618 78102 691174
rect 77546 654618 78102 655174
rect 77546 618618 78102 619174
rect 77546 582618 78102 583174
rect 77546 546618 78102 547174
rect 77546 510618 78102 511174
rect 77546 474618 78102 475174
rect 77546 438618 78102 439174
rect 77546 402618 78102 403174
rect 77546 366618 78102 367174
rect 77546 330618 78102 331174
rect 77546 294618 78102 295174
rect 77546 258618 78102 259174
rect 77546 222618 78102 223174
rect 77546 186618 78102 187174
rect 77546 150618 78102 151174
rect 77546 114618 78102 115174
rect 77546 78618 78102 79174
rect 77546 42618 78102 43174
rect 77546 6618 78102 7174
rect 77546 -2822 78102 -2266
rect 81266 694338 81822 694894
rect 81266 658338 81822 658894
rect 81266 622338 81822 622894
rect 81266 586338 81822 586894
rect 81266 550338 81822 550894
rect 81266 514338 81822 514894
rect 81266 478338 81822 478894
rect 81266 442338 81822 442894
rect 81266 406338 81822 406894
rect 81266 370338 81822 370894
rect 81266 334338 81822 334894
rect 81266 298338 81822 298894
rect 81266 262338 81822 262894
rect 81266 226338 81822 226894
rect 81266 190338 81822 190894
rect 81266 154338 81822 154894
rect 81266 118338 81822 118894
rect 81266 82338 81822 82894
rect 81266 46338 81822 46894
rect 81266 10338 81822 10894
rect 81266 -4742 81822 -4186
rect 102986 711002 103542 711558
rect 99266 709082 99822 709638
rect 95546 707162 96102 707718
rect 84986 698058 85542 698614
rect 84986 662058 85542 662614
rect 84986 626058 85542 626614
rect 84986 590058 85542 590614
rect 84986 554058 85542 554614
rect 84986 518058 85542 518614
rect 84986 482058 85542 482614
rect 84986 446058 85542 446614
rect 84986 410058 85542 410614
rect 84986 374058 85542 374614
rect 84986 338058 85542 338614
rect 84986 302058 85542 302614
rect 84986 266058 85542 266614
rect 84986 230058 85542 230614
rect 84986 194058 85542 194614
rect 84986 158058 85542 158614
rect 84986 122058 85542 122614
rect 84986 86058 85542 86614
rect 84986 50058 85542 50614
rect 84986 14058 85542 14614
rect 66986 -7622 67542 -7066
rect 91826 705242 92382 705798
rect 91826 668898 92382 669454
rect 91826 632898 92382 633454
rect 91826 596898 92382 597454
rect 91826 560898 92382 561454
rect 91826 524898 92382 525454
rect 91826 488898 92382 489454
rect 91826 452898 92382 453454
rect 91826 416898 92382 417454
rect 91826 380898 92382 381454
rect 91826 344898 92382 345454
rect 91826 308898 92382 309454
rect 91826 272898 92382 273454
rect 91826 236898 92382 237454
rect 91826 200898 92382 201454
rect 91826 164898 92382 165454
rect 91826 128898 92382 129454
rect 91826 92898 92382 93454
rect 91826 56898 92382 57454
rect 91826 20898 92382 21454
rect 91826 -1862 92382 -1306
rect 95546 672618 96102 673174
rect 95546 636618 96102 637174
rect 95546 600618 96102 601174
rect 95546 564618 96102 565174
rect 95546 528618 96102 529174
rect 95546 492618 96102 493174
rect 95546 456618 96102 457174
rect 95546 420618 96102 421174
rect 95546 384618 96102 385174
rect 95546 348618 96102 349174
rect 95546 312618 96102 313174
rect 95546 276618 96102 277174
rect 95546 240618 96102 241174
rect 95546 204618 96102 205174
rect 95546 168618 96102 169174
rect 95546 132618 96102 133174
rect 95546 96618 96102 97174
rect 95546 60618 96102 61174
rect 95546 24618 96102 25174
rect 95546 -3782 96102 -3226
rect 99266 676338 99822 676894
rect 99266 640338 99822 640894
rect 99266 604338 99822 604894
rect 99266 568338 99822 568894
rect 99266 532338 99822 532894
rect 99266 496338 99822 496894
rect 99266 460338 99822 460894
rect 99266 424338 99822 424894
rect 99266 388338 99822 388894
rect 99266 352338 99822 352894
rect 99266 316338 99822 316894
rect 99266 280338 99822 280894
rect 99266 244338 99822 244894
rect 99266 208338 99822 208894
rect 99266 172338 99822 172894
rect 99266 136338 99822 136894
rect 99266 100338 99822 100894
rect 99266 64338 99822 64894
rect 99266 28338 99822 28894
rect 99266 -5702 99822 -5146
rect 120986 710042 121542 710598
rect 117266 708122 117822 708678
rect 113546 706202 114102 706758
rect 102986 680058 103542 680614
rect 102986 644058 103542 644614
rect 102986 608058 103542 608614
rect 102986 572058 103542 572614
rect 102986 536058 103542 536614
rect 102986 500058 103542 500614
rect 102986 464058 103542 464614
rect 102986 428058 103542 428614
rect 102986 392058 103542 392614
rect 102986 356058 103542 356614
rect 102986 320058 103542 320614
rect 102986 284058 103542 284614
rect 102986 248058 103542 248614
rect 102986 212058 103542 212614
rect 102986 176058 103542 176614
rect 102986 140058 103542 140614
rect 102986 104058 103542 104614
rect 102986 68058 103542 68614
rect 102986 32058 103542 32614
rect 84986 -6662 85542 -6106
rect 109826 704282 110382 704838
rect 109826 686898 110382 687454
rect 109826 650898 110382 651454
rect 109826 614898 110382 615454
rect 109826 578898 110382 579454
rect 109826 542898 110382 543454
rect 109826 506898 110382 507454
rect 109826 470898 110382 471454
rect 109826 434898 110382 435454
rect 109826 398898 110382 399454
rect 109826 362898 110382 363454
rect 109826 326898 110382 327454
rect 109826 290898 110382 291454
rect 109826 254898 110382 255454
rect 109826 218898 110382 219454
rect 109826 182898 110382 183454
rect 109826 146898 110382 147454
rect 109826 110898 110382 111454
rect 109826 74898 110382 75454
rect 109826 38898 110382 39454
rect 109826 2898 110382 3454
rect 109826 -902 110382 -346
rect 113546 690618 114102 691174
rect 113546 654618 114102 655174
rect 113546 618618 114102 619174
rect 113546 582618 114102 583174
rect 113546 546618 114102 547174
rect 113546 510618 114102 511174
rect 113546 474618 114102 475174
rect 113546 438618 114102 439174
rect 113546 402618 114102 403174
rect 113546 366618 114102 367174
rect 113546 330618 114102 331174
rect 113546 294618 114102 295174
rect 113546 258618 114102 259174
rect 113546 222618 114102 223174
rect 113546 186618 114102 187174
rect 113546 150618 114102 151174
rect 113546 114618 114102 115174
rect 113546 78618 114102 79174
rect 113546 42618 114102 43174
rect 113546 6618 114102 7174
rect 113546 -2822 114102 -2266
rect 117266 694338 117822 694894
rect 117266 658338 117822 658894
rect 117266 622338 117822 622894
rect 117266 586338 117822 586894
rect 117266 550338 117822 550894
rect 117266 514338 117822 514894
rect 117266 478338 117822 478894
rect 117266 442338 117822 442894
rect 117266 406338 117822 406894
rect 117266 370338 117822 370894
rect 117266 334338 117822 334894
rect 117266 298338 117822 298894
rect 117266 262338 117822 262894
rect 117266 226338 117822 226894
rect 117266 190338 117822 190894
rect 117266 154338 117822 154894
rect 117266 118338 117822 118894
rect 117266 82338 117822 82894
rect 117266 46338 117822 46894
rect 117266 10338 117822 10894
rect 117266 -4742 117822 -4186
rect 138986 711002 139542 711558
rect 135266 709082 135822 709638
rect 131546 707162 132102 707718
rect 120986 698058 121542 698614
rect 120986 662058 121542 662614
rect 120986 626058 121542 626614
rect 120986 590058 121542 590614
rect 120986 554058 121542 554614
rect 120986 518058 121542 518614
rect 120986 482058 121542 482614
rect 120986 446058 121542 446614
rect 120986 410058 121542 410614
rect 120986 374058 121542 374614
rect 120986 338058 121542 338614
rect 120986 302058 121542 302614
rect 120986 266058 121542 266614
rect 120986 230058 121542 230614
rect 120986 194058 121542 194614
rect 120986 158058 121542 158614
rect 120986 122058 121542 122614
rect 120986 86058 121542 86614
rect 120986 50058 121542 50614
rect 120986 14058 121542 14614
rect 102986 -7622 103542 -7066
rect 127826 705242 128382 705798
rect 127826 668898 128382 669454
rect 127826 632898 128382 633454
rect 127826 596898 128382 597454
rect 127826 560898 128382 561454
rect 127826 524898 128382 525454
rect 127826 488898 128382 489454
rect 127826 452898 128382 453454
rect 127826 416898 128382 417454
rect 127826 380898 128382 381454
rect 127826 344898 128382 345454
rect 127826 308898 128382 309454
rect 127826 272898 128382 273454
rect 127826 236898 128382 237454
rect 127826 200898 128382 201454
rect 127826 164898 128382 165454
rect 127826 128898 128382 129454
rect 127826 92898 128382 93454
rect 127826 56898 128382 57454
rect 127826 20898 128382 21454
rect 127826 -1862 128382 -1306
rect 131546 672618 132102 673174
rect 131546 636618 132102 637174
rect 131546 600618 132102 601174
rect 131546 564618 132102 565174
rect 131546 528618 132102 529174
rect 131546 492618 132102 493174
rect 131546 456618 132102 457174
rect 131546 420618 132102 421174
rect 131546 384618 132102 385174
rect 131546 348618 132102 349174
rect 131546 312618 132102 313174
rect 131546 276618 132102 277174
rect 131546 240618 132102 241174
rect 131546 204618 132102 205174
rect 131546 168618 132102 169174
rect 131546 132618 132102 133174
rect 131546 96618 132102 97174
rect 131546 60618 132102 61174
rect 131546 24618 132102 25174
rect 131546 -3782 132102 -3226
rect 135266 676338 135822 676894
rect 135266 640338 135822 640894
rect 135266 604338 135822 604894
rect 135266 568338 135822 568894
rect 135266 532338 135822 532894
rect 135266 496338 135822 496894
rect 135266 460338 135822 460894
rect 135266 424338 135822 424894
rect 135266 388338 135822 388894
rect 135266 352338 135822 352894
rect 135266 316338 135822 316894
rect 135266 280338 135822 280894
rect 135266 244338 135822 244894
rect 135266 208338 135822 208894
rect 135266 172338 135822 172894
rect 135266 136338 135822 136894
rect 135266 100338 135822 100894
rect 135266 64338 135822 64894
rect 135266 28338 135822 28894
rect 135266 -5702 135822 -5146
rect 156986 710042 157542 710598
rect 153266 708122 153822 708678
rect 149546 706202 150102 706758
rect 138986 680058 139542 680614
rect 138986 644058 139542 644614
rect 138986 608058 139542 608614
rect 138986 572058 139542 572614
rect 138986 536058 139542 536614
rect 138986 500058 139542 500614
rect 138986 464058 139542 464614
rect 138986 428058 139542 428614
rect 138986 392058 139542 392614
rect 138986 356058 139542 356614
rect 138986 320058 139542 320614
rect 138986 284058 139542 284614
rect 138986 248058 139542 248614
rect 138986 212058 139542 212614
rect 138986 176058 139542 176614
rect 138986 140058 139542 140614
rect 138986 104058 139542 104614
rect 138986 68058 139542 68614
rect 138986 32058 139542 32614
rect 120986 -6662 121542 -6106
rect 145826 704282 146382 704838
rect 145826 686898 146382 687454
rect 145826 650898 146382 651454
rect 145826 614898 146382 615454
rect 145826 578898 146382 579454
rect 145826 542898 146382 543454
rect 145826 506898 146382 507454
rect 145826 470898 146382 471454
rect 145826 434898 146382 435454
rect 145826 398898 146382 399454
rect 145826 362898 146382 363454
rect 145826 326898 146382 327454
rect 145826 290898 146382 291454
rect 145826 254898 146382 255454
rect 145826 218898 146382 219454
rect 145826 182898 146382 183454
rect 145826 146898 146382 147454
rect 145826 110898 146382 111454
rect 145826 74898 146382 75454
rect 145826 38898 146382 39454
rect 145826 2898 146382 3454
rect 145826 -902 146382 -346
rect 149546 690618 150102 691174
rect 149546 654618 150102 655174
rect 149546 618618 150102 619174
rect 149546 582618 150102 583174
rect 149546 546618 150102 547174
rect 149546 510618 150102 511174
rect 149546 474618 150102 475174
rect 149546 438618 150102 439174
rect 149546 402618 150102 403174
rect 149546 366618 150102 367174
rect 149546 330618 150102 331174
rect 149546 294618 150102 295174
rect 149546 258618 150102 259174
rect 149546 222618 150102 223174
rect 149546 186618 150102 187174
rect 149546 150618 150102 151174
rect 149546 114618 150102 115174
rect 149546 78618 150102 79174
rect 149546 42618 150102 43174
rect 149546 6618 150102 7174
rect 149546 -2822 150102 -2266
rect 153266 694338 153822 694894
rect 153266 658338 153822 658894
rect 153266 622338 153822 622894
rect 153266 586338 153822 586894
rect 153266 550338 153822 550894
rect 153266 514338 153822 514894
rect 153266 478338 153822 478894
rect 153266 442338 153822 442894
rect 153266 406338 153822 406894
rect 153266 370338 153822 370894
rect 153266 334338 153822 334894
rect 153266 298338 153822 298894
rect 153266 262338 153822 262894
rect 153266 226338 153822 226894
rect 153266 190338 153822 190894
rect 153266 154338 153822 154894
rect 153266 118338 153822 118894
rect 153266 82338 153822 82894
rect 153266 46338 153822 46894
rect 153266 10338 153822 10894
rect 153266 -4742 153822 -4186
rect 174986 711002 175542 711558
rect 171266 709082 171822 709638
rect 167546 707162 168102 707718
rect 156986 698058 157542 698614
rect 156986 662058 157542 662614
rect 156986 626058 157542 626614
rect 156986 590058 157542 590614
rect 156986 554058 157542 554614
rect 156986 518058 157542 518614
rect 156986 482058 157542 482614
rect 156986 446058 157542 446614
rect 156986 410058 157542 410614
rect 156986 374058 157542 374614
rect 156986 338058 157542 338614
rect 156986 302058 157542 302614
rect 156986 266058 157542 266614
rect 156986 230058 157542 230614
rect 156986 194058 157542 194614
rect 156986 158058 157542 158614
rect 156986 122058 157542 122614
rect 156986 86058 157542 86614
rect 156986 50058 157542 50614
rect 156986 14058 157542 14614
rect 138986 -7622 139542 -7066
rect 163826 705242 164382 705798
rect 163826 668898 164382 669454
rect 163826 632898 164382 633454
rect 163826 596898 164382 597454
rect 163826 560898 164382 561454
rect 163826 524898 164382 525454
rect 163826 488898 164382 489454
rect 163826 452898 164382 453454
rect 163826 416898 164382 417454
rect 163826 380898 164382 381454
rect 163826 344898 164382 345454
rect 163826 308898 164382 309454
rect 163826 272898 164382 273454
rect 163826 236898 164382 237454
rect 163826 200898 164382 201454
rect 163826 164898 164382 165454
rect 163826 128898 164382 129454
rect 163826 92898 164382 93454
rect 163826 56898 164382 57454
rect 163826 20898 164382 21454
rect 163826 -1862 164382 -1306
rect 167546 672618 168102 673174
rect 167546 636618 168102 637174
rect 167546 600618 168102 601174
rect 167546 564618 168102 565174
rect 167546 528618 168102 529174
rect 167546 492618 168102 493174
rect 167546 456618 168102 457174
rect 167546 420618 168102 421174
rect 167546 384618 168102 385174
rect 167546 348618 168102 349174
rect 167546 312618 168102 313174
rect 167546 276618 168102 277174
rect 167546 240618 168102 241174
rect 167546 204618 168102 205174
rect 167546 168618 168102 169174
rect 167546 132618 168102 133174
rect 167546 96618 168102 97174
rect 167546 60618 168102 61174
rect 167546 24618 168102 25174
rect 167546 -3782 168102 -3226
rect 171266 676338 171822 676894
rect 171266 640338 171822 640894
rect 171266 604338 171822 604894
rect 171266 568338 171822 568894
rect 171266 532338 171822 532894
rect 171266 496338 171822 496894
rect 171266 460338 171822 460894
rect 171266 424338 171822 424894
rect 171266 388338 171822 388894
rect 171266 352338 171822 352894
rect 171266 316338 171822 316894
rect 171266 280338 171822 280894
rect 171266 244338 171822 244894
rect 171266 208338 171822 208894
rect 171266 172338 171822 172894
rect 171266 136338 171822 136894
rect 171266 100338 171822 100894
rect 171266 64338 171822 64894
rect 171266 28338 171822 28894
rect 171266 -5702 171822 -5146
rect 192986 710042 193542 710598
rect 189266 708122 189822 708678
rect 185546 706202 186102 706758
rect 174986 680058 175542 680614
rect 174986 644058 175542 644614
rect 174986 608058 175542 608614
rect 174986 572058 175542 572614
rect 174986 536058 175542 536614
rect 174986 500058 175542 500614
rect 174986 464058 175542 464614
rect 174986 428058 175542 428614
rect 174986 392058 175542 392614
rect 174986 356058 175542 356614
rect 174986 320058 175542 320614
rect 174986 284058 175542 284614
rect 174986 248058 175542 248614
rect 174986 212058 175542 212614
rect 174986 176058 175542 176614
rect 174986 140058 175542 140614
rect 174986 104058 175542 104614
rect 174986 68058 175542 68614
rect 174986 32058 175542 32614
rect 156986 -6662 157542 -6106
rect 181826 704282 182382 704838
rect 181826 686898 182382 687454
rect 181826 650898 182382 651454
rect 181826 614898 182382 615454
rect 181826 578898 182382 579454
rect 181826 542898 182382 543454
rect 181826 506898 182382 507454
rect 181826 470898 182382 471454
rect 181826 434898 182382 435454
rect 181826 398898 182382 399454
rect 181826 362898 182382 363454
rect 181826 326898 182382 327454
rect 181826 290898 182382 291454
rect 181826 254898 182382 255454
rect 181826 218898 182382 219454
rect 181826 182898 182382 183454
rect 181826 146898 182382 147454
rect 181826 110898 182382 111454
rect 181826 74898 182382 75454
rect 181826 38898 182382 39454
rect 181826 2898 182382 3454
rect 181826 -902 182382 -346
rect 185546 690618 186102 691174
rect 185546 654618 186102 655174
rect 185546 618618 186102 619174
rect 185546 582618 186102 583174
rect 185546 546618 186102 547174
rect 185546 510618 186102 511174
rect 185546 474618 186102 475174
rect 185546 438618 186102 439174
rect 185546 402618 186102 403174
rect 185546 366618 186102 367174
rect 185546 330618 186102 331174
rect 185546 294618 186102 295174
rect 185546 258618 186102 259174
rect 185546 222618 186102 223174
rect 185546 186618 186102 187174
rect 185546 150618 186102 151174
rect 185546 114618 186102 115174
rect 185546 78618 186102 79174
rect 185546 42618 186102 43174
rect 185546 6618 186102 7174
rect 185546 -2822 186102 -2266
rect 189266 694338 189822 694894
rect 189266 658338 189822 658894
rect 189266 622338 189822 622894
rect 189266 586338 189822 586894
rect 189266 550338 189822 550894
rect 189266 514338 189822 514894
rect 189266 478338 189822 478894
rect 189266 442338 189822 442894
rect 189266 406338 189822 406894
rect 189266 370338 189822 370894
rect 189266 334338 189822 334894
rect 189266 298338 189822 298894
rect 189266 262338 189822 262894
rect 189266 226338 189822 226894
rect 189266 190338 189822 190894
rect 189266 154338 189822 154894
rect 189266 118338 189822 118894
rect 189266 82338 189822 82894
rect 189266 46338 189822 46894
rect 189266 10338 189822 10894
rect 189266 -4742 189822 -4186
rect 210986 711002 211542 711558
rect 207266 709082 207822 709638
rect 203546 707162 204102 707718
rect 192986 698058 193542 698614
rect 192986 662058 193542 662614
rect 192986 626058 193542 626614
rect 192986 590058 193542 590614
rect 192986 554058 193542 554614
rect 192986 518058 193542 518614
rect 192986 482058 193542 482614
rect 192986 446058 193542 446614
rect 192986 410058 193542 410614
rect 192986 374058 193542 374614
rect 192986 338058 193542 338614
rect 192986 302058 193542 302614
rect 192986 266058 193542 266614
rect 192986 230058 193542 230614
rect 192986 194058 193542 194614
rect 192986 158058 193542 158614
rect 192986 122058 193542 122614
rect 192986 86058 193542 86614
rect 192986 50058 193542 50614
rect 192986 14058 193542 14614
rect 174986 -7622 175542 -7066
rect 199826 705242 200382 705798
rect 199826 668898 200382 669454
rect 199826 632898 200382 633454
rect 199826 596898 200382 597454
rect 199826 560898 200382 561454
rect 199826 524898 200382 525454
rect 199826 488898 200382 489454
rect 199826 452898 200382 453454
rect 199826 416898 200382 417454
rect 199826 380898 200382 381454
rect 199826 344898 200382 345454
rect 199826 308898 200382 309454
rect 199826 272898 200382 273454
rect 199826 236898 200382 237454
rect 199826 200898 200382 201454
rect 199826 164898 200382 165454
rect 199826 128898 200382 129454
rect 199826 92898 200382 93454
rect 199826 56898 200382 57454
rect 199826 20898 200382 21454
rect 199826 -1862 200382 -1306
rect 203546 672618 204102 673174
rect 203546 636618 204102 637174
rect 203546 600618 204102 601174
rect 203546 564618 204102 565174
rect 203546 528618 204102 529174
rect 203546 492618 204102 493174
rect 203546 456618 204102 457174
rect 203546 420618 204102 421174
rect 203546 384618 204102 385174
rect 203546 348618 204102 349174
rect 203546 312618 204102 313174
rect 203546 276618 204102 277174
rect 203546 240618 204102 241174
rect 203546 204618 204102 205174
rect 203546 168618 204102 169174
rect 203546 132618 204102 133174
rect 203546 96618 204102 97174
rect 203546 60618 204102 61174
rect 203546 24618 204102 25174
rect 203546 -3782 204102 -3226
rect 207266 676338 207822 676894
rect 207266 640338 207822 640894
rect 207266 604338 207822 604894
rect 207266 568338 207822 568894
rect 207266 532338 207822 532894
rect 207266 496338 207822 496894
rect 207266 460338 207822 460894
rect 207266 424338 207822 424894
rect 207266 388338 207822 388894
rect 207266 352338 207822 352894
rect 207266 316338 207822 316894
rect 207266 280338 207822 280894
rect 207266 244338 207822 244894
rect 207266 208338 207822 208894
rect 207266 172338 207822 172894
rect 207266 136338 207822 136894
rect 207266 100338 207822 100894
rect 207266 64338 207822 64894
rect 207266 28338 207822 28894
rect 207266 -5702 207822 -5146
rect 228986 710042 229542 710598
rect 225266 708122 225822 708678
rect 221546 706202 222102 706758
rect 210986 680058 211542 680614
rect 210986 644058 211542 644614
rect 210986 608058 211542 608614
rect 210986 572058 211542 572614
rect 210986 536058 211542 536614
rect 210986 500058 211542 500614
rect 210986 464058 211542 464614
rect 210986 428058 211542 428614
rect 210986 392058 211542 392614
rect 210986 356058 211542 356614
rect 210986 320058 211542 320614
rect 210986 284058 211542 284614
rect 210986 248058 211542 248614
rect 210986 212058 211542 212614
rect 210986 176058 211542 176614
rect 210986 140058 211542 140614
rect 210986 104058 211542 104614
rect 210986 68058 211542 68614
rect 210986 32058 211542 32614
rect 192986 -6662 193542 -6106
rect 217826 704282 218382 704838
rect 217826 686898 218382 687454
rect 217826 650898 218382 651454
rect 217826 614898 218382 615454
rect 217826 578898 218382 579454
rect 217826 542898 218382 543454
rect 217826 506898 218382 507454
rect 217826 470898 218382 471454
rect 217826 434898 218382 435454
rect 217826 398898 218382 399454
rect 217826 362898 218382 363454
rect 217826 326898 218382 327454
rect 217826 290898 218382 291454
rect 217826 254898 218382 255454
rect 217826 218898 218382 219454
rect 217826 182898 218382 183454
rect 217826 146898 218382 147454
rect 217826 110898 218382 111454
rect 217826 74898 218382 75454
rect 217826 38898 218382 39454
rect 217826 2898 218382 3454
rect 217826 -902 218382 -346
rect 221546 690618 222102 691174
rect 221546 654618 222102 655174
rect 221546 618618 222102 619174
rect 221546 582618 222102 583174
rect 221546 546618 222102 547174
rect 221546 510618 222102 511174
rect 221546 474618 222102 475174
rect 221546 438618 222102 439174
rect 221546 402618 222102 403174
rect 221546 366618 222102 367174
rect 221546 330618 222102 331174
rect 221546 294618 222102 295174
rect 221546 258618 222102 259174
rect 221546 222618 222102 223174
rect 221546 186618 222102 187174
rect 221546 150618 222102 151174
rect 221546 114618 222102 115174
rect 221546 78618 222102 79174
rect 221546 42618 222102 43174
rect 221546 6618 222102 7174
rect 221546 -2822 222102 -2266
rect 225266 694338 225822 694894
rect 225266 658338 225822 658894
rect 225266 622338 225822 622894
rect 225266 586338 225822 586894
rect 225266 550338 225822 550894
rect 225266 514338 225822 514894
rect 225266 478338 225822 478894
rect 225266 442338 225822 442894
rect 225266 406338 225822 406894
rect 225266 370338 225822 370894
rect 225266 334338 225822 334894
rect 225266 298338 225822 298894
rect 225266 262338 225822 262894
rect 225266 226338 225822 226894
rect 225266 190338 225822 190894
rect 225266 154338 225822 154894
rect 225266 118338 225822 118894
rect 225266 82338 225822 82894
rect 225266 46338 225822 46894
rect 225266 10338 225822 10894
rect 225266 -4742 225822 -4186
rect 246986 711002 247542 711558
rect 243266 709082 243822 709638
rect 239546 707162 240102 707718
rect 228986 698058 229542 698614
rect 228986 662058 229542 662614
rect 228986 626058 229542 626614
rect 228986 590058 229542 590614
rect 228986 554058 229542 554614
rect 228986 518058 229542 518614
rect 228986 482058 229542 482614
rect 235826 705242 236382 705798
rect 235826 668898 236382 669454
rect 235826 632898 236382 633454
rect 235826 596898 236382 597454
rect 235826 560898 236382 561454
rect 235826 524898 236382 525454
rect 235826 488898 236382 489454
rect 239546 672618 240102 673174
rect 239546 636618 240102 637174
rect 239546 600618 240102 601174
rect 239546 564618 240102 565174
rect 239546 528618 240102 529174
rect 239546 492618 240102 493174
rect 243266 676338 243822 676894
rect 243266 640338 243822 640894
rect 243266 604338 243822 604894
rect 243266 568338 243822 568894
rect 243266 532338 243822 532894
rect 243266 496338 243822 496894
rect 243266 460338 243822 460894
rect 264986 710042 265542 710598
rect 261266 708122 261822 708678
rect 257546 706202 258102 706758
rect 246986 680058 247542 680614
rect 246986 644058 247542 644614
rect 246986 608058 247542 608614
rect 246986 572058 247542 572614
rect 246986 536058 247542 536614
rect 246986 500058 247542 500614
rect 246986 464058 247542 464614
rect 253826 704282 254382 704838
rect 253826 686898 254382 687454
rect 253826 650898 254382 651454
rect 253826 614898 254382 615454
rect 253826 578898 254382 579454
rect 253826 542898 254382 543454
rect 253826 506898 254382 507454
rect 253826 470898 254382 471454
rect 257546 690618 258102 691174
rect 257546 654618 258102 655174
rect 257546 618618 258102 619174
rect 257546 582618 258102 583174
rect 257546 546618 258102 547174
rect 257546 510618 258102 511174
rect 257546 474618 258102 475174
rect 261266 694338 261822 694894
rect 261266 658338 261822 658894
rect 261266 622338 261822 622894
rect 261266 586338 261822 586894
rect 261266 550338 261822 550894
rect 261266 514338 261822 514894
rect 261266 478338 261822 478894
rect 282986 711002 283542 711558
rect 279266 709082 279822 709638
rect 275546 707162 276102 707718
rect 264986 698058 265542 698614
rect 264986 662058 265542 662614
rect 264986 626058 265542 626614
rect 264986 590058 265542 590614
rect 264986 554058 265542 554614
rect 264986 518058 265542 518614
rect 264986 482058 265542 482614
rect 271826 705242 272382 705798
rect 271826 668898 272382 669454
rect 271826 632898 272382 633454
rect 271826 596898 272382 597454
rect 271826 560898 272382 561454
rect 271826 524898 272382 525454
rect 271826 488898 272382 489454
rect 275546 672618 276102 673174
rect 275546 636618 276102 637174
rect 275546 600618 276102 601174
rect 275546 564618 276102 565174
rect 275546 528618 276102 529174
rect 275546 492618 276102 493174
rect 279266 676338 279822 676894
rect 279266 640338 279822 640894
rect 279266 604338 279822 604894
rect 279266 568338 279822 568894
rect 279266 532338 279822 532894
rect 279266 496338 279822 496894
rect 279266 460338 279822 460894
rect 300986 710042 301542 710598
rect 297266 708122 297822 708678
rect 293546 706202 294102 706758
rect 282986 680058 283542 680614
rect 282986 644058 283542 644614
rect 282986 608058 283542 608614
rect 282986 572058 283542 572614
rect 282986 536058 283542 536614
rect 282986 500058 283542 500614
rect 282986 464058 283542 464614
rect 289826 704282 290382 704838
rect 289826 686898 290382 687454
rect 289826 650898 290382 651454
rect 289826 614898 290382 615454
rect 289826 578898 290382 579454
rect 289826 542898 290382 543454
rect 289826 506898 290382 507454
rect 289826 470898 290382 471454
rect 293546 690618 294102 691174
rect 293546 654618 294102 655174
rect 293546 618618 294102 619174
rect 293546 582618 294102 583174
rect 293546 546618 294102 547174
rect 293546 510618 294102 511174
rect 293546 474618 294102 475174
rect 297266 694338 297822 694894
rect 297266 658338 297822 658894
rect 297266 622338 297822 622894
rect 297266 586338 297822 586894
rect 297266 550338 297822 550894
rect 297266 514338 297822 514894
rect 297266 478338 297822 478894
rect 318986 711002 319542 711558
rect 315266 709082 315822 709638
rect 311546 707162 312102 707718
rect 300986 698058 301542 698614
rect 300986 662058 301542 662614
rect 300986 626058 301542 626614
rect 300986 590058 301542 590614
rect 300986 554058 301542 554614
rect 300986 518058 301542 518614
rect 300986 482058 301542 482614
rect 307826 705242 308382 705798
rect 307826 668898 308382 669454
rect 307826 632898 308382 633454
rect 307826 596898 308382 597454
rect 307826 560898 308382 561454
rect 307826 524898 308382 525454
rect 307826 488898 308382 489454
rect 311546 672618 312102 673174
rect 311546 636618 312102 637174
rect 311546 600618 312102 601174
rect 311546 564618 312102 565174
rect 311546 528618 312102 529174
rect 311546 492618 312102 493174
rect 315266 676338 315822 676894
rect 315266 640338 315822 640894
rect 315266 604338 315822 604894
rect 315266 568338 315822 568894
rect 315266 532338 315822 532894
rect 315266 496338 315822 496894
rect 315266 460338 315822 460894
rect 336986 710042 337542 710598
rect 333266 708122 333822 708678
rect 329546 706202 330102 706758
rect 318986 680058 319542 680614
rect 318986 644058 319542 644614
rect 318986 608058 319542 608614
rect 318986 572058 319542 572614
rect 318986 536058 319542 536614
rect 318986 500058 319542 500614
rect 318986 464058 319542 464614
rect 325826 704282 326382 704838
rect 325826 686898 326382 687454
rect 325826 650898 326382 651454
rect 325826 614898 326382 615454
rect 325826 578898 326382 579454
rect 325826 542898 326382 543454
rect 325826 506898 326382 507454
rect 325826 470898 326382 471454
rect 329546 690618 330102 691174
rect 329546 654618 330102 655174
rect 329546 618618 330102 619174
rect 329546 582618 330102 583174
rect 329546 546618 330102 547174
rect 329546 510618 330102 511174
rect 329546 474618 330102 475174
rect 333266 694338 333822 694894
rect 333266 658338 333822 658894
rect 333266 622338 333822 622894
rect 333266 586338 333822 586894
rect 333266 550338 333822 550894
rect 333266 514338 333822 514894
rect 333266 478338 333822 478894
rect 354986 711002 355542 711558
rect 351266 709082 351822 709638
rect 347546 707162 348102 707718
rect 336986 698058 337542 698614
rect 336986 662058 337542 662614
rect 336986 626058 337542 626614
rect 336986 590058 337542 590614
rect 336986 554058 337542 554614
rect 336986 518058 337542 518614
rect 336986 482058 337542 482614
rect 343826 705242 344382 705798
rect 343826 668898 344382 669454
rect 343826 632898 344382 633454
rect 343826 596898 344382 597454
rect 343826 560898 344382 561454
rect 343826 524898 344382 525454
rect 343826 488898 344382 489454
rect 347546 672618 348102 673174
rect 347546 636618 348102 637174
rect 347546 600618 348102 601174
rect 347546 564618 348102 565174
rect 347546 528618 348102 529174
rect 347546 492618 348102 493174
rect 351266 676338 351822 676894
rect 351266 640338 351822 640894
rect 351266 604338 351822 604894
rect 351266 568338 351822 568894
rect 351266 532338 351822 532894
rect 351266 496338 351822 496894
rect 351266 460338 351822 460894
rect 372986 710042 373542 710598
rect 369266 708122 369822 708678
rect 365546 706202 366102 706758
rect 354986 680058 355542 680614
rect 354986 644058 355542 644614
rect 354986 608058 355542 608614
rect 354986 572058 355542 572614
rect 354986 536058 355542 536614
rect 354986 500058 355542 500614
rect 354986 464058 355542 464614
rect 361826 704282 362382 704838
rect 361826 686898 362382 687454
rect 361826 650898 362382 651454
rect 361826 614898 362382 615454
rect 361826 578898 362382 579454
rect 361826 542898 362382 543454
rect 361826 506898 362382 507454
rect 361826 470898 362382 471454
rect 365546 690618 366102 691174
rect 365546 654618 366102 655174
rect 365546 618618 366102 619174
rect 365546 582618 366102 583174
rect 365546 546618 366102 547174
rect 365546 510618 366102 511174
rect 365546 474618 366102 475174
rect 369266 694338 369822 694894
rect 369266 658338 369822 658894
rect 369266 622338 369822 622894
rect 369266 586338 369822 586894
rect 369266 550338 369822 550894
rect 369266 514338 369822 514894
rect 369266 478338 369822 478894
rect 390986 711002 391542 711558
rect 387266 709082 387822 709638
rect 383546 707162 384102 707718
rect 372986 698058 373542 698614
rect 372986 662058 373542 662614
rect 372986 626058 373542 626614
rect 372986 590058 373542 590614
rect 372986 554058 373542 554614
rect 372986 518058 373542 518614
rect 372986 482058 373542 482614
rect 379826 705242 380382 705798
rect 379826 668898 380382 669454
rect 379826 632898 380382 633454
rect 379826 596898 380382 597454
rect 379826 560898 380382 561454
rect 379826 524898 380382 525454
rect 379826 488898 380382 489454
rect 383546 672618 384102 673174
rect 383546 636618 384102 637174
rect 383546 600618 384102 601174
rect 383546 564618 384102 565174
rect 383546 528618 384102 529174
rect 383546 492618 384102 493174
rect 387266 676338 387822 676894
rect 387266 640338 387822 640894
rect 387266 604338 387822 604894
rect 387266 568338 387822 568894
rect 387266 532338 387822 532894
rect 387266 496338 387822 496894
rect 387266 460338 387822 460894
rect 408986 710042 409542 710598
rect 405266 708122 405822 708678
rect 401546 706202 402102 706758
rect 390986 680058 391542 680614
rect 390986 644058 391542 644614
rect 390986 608058 391542 608614
rect 390986 572058 391542 572614
rect 390986 536058 391542 536614
rect 390986 500058 391542 500614
rect 390986 464058 391542 464614
rect 397826 704282 398382 704838
rect 397826 686898 398382 687454
rect 397826 650898 398382 651454
rect 397826 614898 398382 615454
rect 397826 578898 398382 579454
rect 397826 542898 398382 543454
rect 397826 506898 398382 507454
rect 397826 470898 398382 471454
rect 401546 690618 402102 691174
rect 401546 654618 402102 655174
rect 401546 618618 402102 619174
rect 401546 582618 402102 583174
rect 401546 546618 402102 547174
rect 401546 510618 402102 511174
rect 401546 474618 402102 475174
rect 405266 694338 405822 694894
rect 405266 658338 405822 658894
rect 405266 622338 405822 622894
rect 405266 586338 405822 586894
rect 405266 550338 405822 550894
rect 405266 514338 405822 514894
rect 405266 478338 405822 478894
rect 426986 711002 427542 711558
rect 423266 709082 423822 709638
rect 419546 707162 420102 707718
rect 408986 698058 409542 698614
rect 408986 662058 409542 662614
rect 408986 626058 409542 626614
rect 408986 590058 409542 590614
rect 408986 554058 409542 554614
rect 408986 518058 409542 518614
rect 408986 482058 409542 482614
rect 415826 705242 416382 705798
rect 415826 668898 416382 669454
rect 415826 632898 416382 633454
rect 415826 596898 416382 597454
rect 415826 560898 416382 561454
rect 415826 524898 416382 525454
rect 415826 488898 416382 489454
rect 228986 446058 229542 446614
rect 228986 410058 229542 410614
rect 228986 374058 229542 374614
rect 228986 338058 229542 338614
rect 228986 302058 229542 302614
rect 228986 266058 229542 266614
rect 228986 230058 229542 230614
rect 228986 194058 229542 194614
rect 228986 158058 229542 158614
rect 228986 122058 229542 122614
rect 228986 86058 229542 86614
rect 228986 50058 229542 50614
rect 228986 14058 229542 14614
rect 210986 -7622 211542 -7066
rect 235826 308898 236382 309454
rect 235826 272898 236382 273454
rect 235826 236898 236382 237454
rect 235826 200898 236382 201454
rect 235826 164898 236382 165454
rect 235826 128898 236382 129454
rect 235826 92898 236382 93454
rect 235826 56898 236382 57454
rect 239250 435218 239486 435454
rect 239250 434898 239486 435134
rect 239250 399218 239486 399454
rect 239250 398898 239486 399134
rect 239250 363218 239486 363454
rect 239250 362898 239486 363134
rect 239546 312618 240102 313174
rect 239546 276618 240102 277174
rect 239546 240618 240102 241174
rect 239546 204618 240102 205174
rect 239546 168618 240102 169174
rect 239546 132618 240102 133174
rect 239546 96618 240102 97174
rect 239546 60618 240102 61174
rect 235826 20898 236382 21454
rect 235826 -1862 236382 -1306
rect 243266 316338 243822 316894
rect 243266 280338 243822 280894
rect 243266 244338 243822 244894
rect 243266 208338 243822 208894
rect 243266 172338 243822 172894
rect 243266 136338 243822 136894
rect 243266 100338 243822 100894
rect 243266 64338 243822 64894
rect 239546 24618 240102 25174
rect 239546 -3782 240102 -3226
rect 246986 320058 247542 320614
rect 246986 284058 247542 284614
rect 246986 248058 247542 248614
rect 246986 212058 247542 212614
rect 246986 176058 247542 176614
rect 246986 140058 247542 140614
rect 246986 104058 247542 104614
rect 254610 453218 254846 453454
rect 254610 452898 254846 453134
rect 254610 417218 254846 417454
rect 254610 416898 254846 417134
rect 254610 381218 254846 381454
rect 254610 380898 254846 381134
rect 254610 345218 254846 345454
rect 254610 344898 254846 345134
rect 253826 326898 254382 327454
rect 253826 290898 254382 291454
rect 253826 254898 254382 255454
rect 253826 218898 254382 219454
rect 253826 182898 254382 183454
rect 257546 330618 258102 331174
rect 257546 294618 258102 295174
rect 257546 258618 258102 259174
rect 257546 222618 258102 223174
rect 261266 334338 261822 334894
rect 261266 298338 261822 298894
rect 261266 262338 261822 262894
rect 261266 226338 261822 226894
rect 257546 186618 258102 187174
rect 253826 146898 254382 147454
rect 253826 110898 254382 111454
rect 246986 68058 247542 68614
rect 243266 28338 243822 28894
rect 243266 -5702 243822 -5146
rect 246986 32058 247542 32614
rect 228986 -6662 229542 -6106
rect 253826 74898 254382 75454
rect 253826 38898 254382 39454
rect 253826 2898 254382 3454
rect 253826 -902 254382 -346
rect 257546 150618 258102 151174
rect 257546 114618 258102 115174
rect 257546 78618 258102 79174
rect 257546 42618 258102 43174
rect 257546 6618 258102 7174
rect 257546 -2822 258102 -2266
rect 264986 302058 265542 302614
rect 264986 266058 265542 266614
rect 285330 453218 285566 453454
rect 285330 452898 285566 453134
rect 316050 453218 316286 453454
rect 316050 452898 316286 453134
rect 346770 453218 347006 453454
rect 346770 452898 347006 453134
rect 377490 453218 377726 453454
rect 377490 452898 377726 453134
rect 269970 435218 270206 435454
rect 269970 434898 270206 435134
rect 300690 435218 300926 435454
rect 300690 434898 300926 435134
rect 331410 435218 331646 435454
rect 331410 434898 331646 435134
rect 362130 435218 362366 435454
rect 362130 434898 362366 435134
rect 285330 417218 285566 417454
rect 285330 416898 285566 417134
rect 316050 417218 316286 417454
rect 316050 416898 316286 417134
rect 346770 417218 347006 417454
rect 346770 416898 347006 417134
rect 377490 417218 377726 417454
rect 377490 416898 377726 417134
rect 269970 399218 270206 399454
rect 269970 398898 270206 399134
rect 300690 399218 300926 399454
rect 300690 398898 300926 399134
rect 331410 399218 331646 399454
rect 331410 398898 331646 399134
rect 362130 399218 362366 399454
rect 362130 398898 362366 399134
rect 285330 381218 285566 381454
rect 285330 380898 285566 381134
rect 316050 381218 316286 381454
rect 316050 380898 316286 381134
rect 346770 381218 347006 381454
rect 346770 380898 347006 381134
rect 377490 381218 377726 381454
rect 377490 380898 377726 381134
rect 269970 363218 270206 363454
rect 269970 362898 270206 363134
rect 300690 363218 300926 363454
rect 300690 362898 300926 363134
rect 331410 363218 331646 363454
rect 331410 362898 331646 363134
rect 362130 363218 362366 363454
rect 362130 362898 362366 363134
rect 285330 345218 285566 345454
rect 285330 344898 285566 345134
rect 316050 345218 316286 345454
rect 316050 344898 316286 345134
rect 346770 345218 347006 345454
rect 346770 344898 347006 345134
rect 377490 345218 377726 345454
rect 377490 344898 377726 345134
rect 271826 308898 272382 309454
rect 271826 272898 272382 273454
rect 264986 230058 265542 230614
rect 261266 190338 261822 190894
rect 261266 154338 261822 154894
rect 261266 118338 261822 118894
rect 261266 82338 261822 82894
rect 261266 46338 261822 46894
rect 261266 10338 261822 10894
rect 261266 -4742 261822 -4186
rect 264986 194058 265542 194614
rect 264986 158058 265542 158614
rect 264986 122058 265542 122614
rect 264986 86058 265542 86614
rect 264986 50058 265542 50614
rect 264986 14058 265542 14614
rect 246986 -7622 247542 -7066
rect 271826 236898 272382 237454
rect 271826 200898 272382 201454
rect 271826 164898 272382 165454
rect 271826 128898 272382 129454
rect 271826 92898 272382 93454
rect 271826 56898 272382 57454
rect 271826 20898 272382 21454
rect 271826 -1862 272382 -1306
rect 275546 312618 276102 313174
rect 275546 276618 276102 277174
rect 275546 240618 276102 241174
rect 275546 204618 276102 205174
rect 275546 168618 276102 169174
rect 275546 132618 276102 133174
rect 275546 96618 276102 97174
rect 275546 60618 276102 61174
rect 275546 24618 276102 25174
rect 275546 -3782 276102 -3226
rect 279266 316338 279822 316894
rect 279266 280338 279822 280894
rect 279266 244338 279822 244894
rect 279266 208338 279822 208894
rect 279266 172338 279822 172894
rect 279266 136338 279822 136894
rect 279266 100338 279822 100894
rect 279266 64338 279822 64894
rect 279266 28338 279822 28894
rect 279266 -5702 279822 -5146
rect 282986 320058 283542 320614
rect 282986 284058 283542 284614
rect 282986 248058 283542 248614
rect 282986 212058 283542 212614
rect 282986 176058 283542 176614
rect 282986 140058 283542 140614
rect 282986 104058 283542 104614
rect 282986 68058 283542 68614
rect 282986 32058 283542 32614
rect 264986 -6662 265542 -6106
rect 289826 326898 290382 327454
rect 289826 290898 290382 291454
rect 289826 254898 290382 255454
rect 289826 218898 290382 219454
rect 289826 182898 290382 183454
rect 289826 146898 290382 147454
rect 289826 110898 290382 111454
rect 289826 74898 290382 75454
rect 289826 38898 290382 39454
rect 289826 2898 290382 3454
rect 289826 -902 290382 -346
rect 293546 330618 294102 331174
rect 293546 294618 294102 295174
rect 293546 258618 294102 259174
rect 293546 222618 294102 223174
rect 293546 186618 294102 187174
rect 293546 150618 294102 151174
rect 293546 114618 294102 115174
rect 293546 78618 294102 79174
rect 293546 42618 294102 43174
rect 293546 6618 294102 7174
rect 293546 -2822 294102 -2266
rect 297266 334338 297822 334894
rect 297266 298338 297822 298894
rect 297266 262338 297822 262894
rect 297266 226338 297822 226894
rect 297266 190338 297822 190894
rect 297266 154338 297822 154894
rect 297266 118338 297822 118894
rect 297266 82338 297822 82894
rect 297266 46338 297822 46894
rect 297266 10338 297822 10894
rect 297266 -4742 297822 -4186
rect 300986 302058 301542 302614
rect 300986 266058 301542 266614
rect 300986 230058 301542 230614
rect 300986 194058 301542 194614
rect 300986 158058 301542 158614
rect 300986 122058 301542 122614
rect 300986 86058 301542 86614
rect 300986 50058 301542 50614
rect 300986 14058 301542 14614
rect 282986 -7622 283542 -7066
rect 307826 308898 308382 309454
rect 307826 272898 308382 273454
rect 307826 236898 308382 237454
rect 307826 200898 308382 201454
rect 307826 164898 308382 165454
rect 307826 128898 308382 129454
rect 307826 92898 308382 93454
rect 307826 56898 308382 57454
rect 307826 20898 308382 21454
rect 307826 -1862 308382 -1306
rect 311546 312618 312102 313174
rect 311546 276618 312102 277174
rect 311546 240618 312102 241174
rect 311546 204618 312102 205174
rect 311546 168618 312102 169174
rect 311546 132618 312102 133174
rect 311546 96618 312102 97174
rect 311546 60618 312102 61174
rect 311546 24618 312102 25174
rect 311546 -3782 312102 -3226
rect 315266 316338 315822 316894
rect 315266 280338 315822 280894
rect 315266 244338 315822 244894
rect 315266 208338 315822 208894
rect 315266 172338 315822 172894
rect 315266 136338 315822 136894
rect 315266 100338 315822 100894
rect 315266 64338 315822 64894
rect 315266 28338 315822 28894
rect 315266 -5702 315822 -5146
rect 318986 320058 319542 320614
rect 318986 284058 319542 284614
rect 318986 248058 319542 248614
rect 318986 212058 319542 212614
rect 318986 176058 319542 176614
rect 318986 140058 319542 140614
rect 318986 104058 319542 104614
rect 318986 68058 319542 68614
rect 318986 32058 319542 32614
rect 300986 -6662 301542 -6106
rect 325826 326898 326382 327454
rect 325826 290898 326382 291454
rect 325826 254898 326382 255454
rect 325826 218898 326382 219454
rect 325826 182898 326382 183454
rect 325826 146898 326382 147454
rect 325826 110898 326382 111454
rect 325826 74898 326382 75454
rect 325826 38898 326382 39454
rect 325826 2898 326382 3454
rect 325826 -902 326382 -346
rect 329546 330618 330102 331174
rect 329546 294618 330102 295174
rect 329546 258618 330102 259174
rect 329546 222618 330102 223174
rect 329546 186618 330102 187174
rect 329546 150618 330102 151174
rect 329546 114618 330102 115174
rect 329546 78618 330102 79174
rect 329546 42618 330102 43174
rect 329546 6618 330102 7174
rect 329546 -2822 330102 -2266
rect 333266 334338 333822 334894
rect 333266 298338 333822 298894
rect 333266 262338 333822 262894
rect 333266 226338 333822 226894
rect 333266 190338 333822 190894
rect 333266 154338 333822 154894
rect 333266 118338 333822 118894
rect 333266 82338 333822 82894
rect 333266 46338 333822 46894
rect 333266 10338 333822 10894
rect 333266 -4742 333822 -4186
rect 336986 302058 337542 302614
rect 336986 266058 337542 266614
rect 336986 230058 337542 230614
rect 336986 194058 337542 194614
rect 336986 158058 337542 158614
rect 336986 122058 337542 122614
rect 336986 86058 337542 86614
rect 336986 50058 337542 50614
rect 336986 14058 337542 14614
rect 318986 -7622 319542 -7066
rect 343826 308898 344382 309454
rect 343826 272898 344382 273454
rect 343826 236898 344382 237454
rect 343826 200898 344382 201454
rect 343826 164898 344382 165454
rect 343826 128898 344382 129454
rect 343826 92898 344382 93454
rect 343826 56898 344382 57454
rect 343826 20898 344382 21454
rect 343826 -1862 344382 -1306
rect 347546 312618 348102 313174
rect 347546 276618 348102 277174
rect 347546 240618 348102 241174
rect 347546 204618 348102 205174
rect 347546 168618 348102 169174
rect 347546 132618 348102 133174
rect 347546 96618 348102 97174
rect 347546 60618 348102 61174
rect 347546 24618 348102 25174
rect 347546 -3782 348102 -3226
rect 351266 316338 351822 316894
rect 351266 280338 351822 280894
rect 351266 244338 351822 244894
rect 351266 208338 351822 208894
rect 351266 172338 351822 172894
rect 351266 136338 351822 136894
rect 351266 100338 351822 100894
rect 351266 64338 351822 64894
rect 351266 28338 351822 28894
rect 351266 -5702 351822 -5146
rect 354986 320058 355542 320614
rect 354986 284058 355542 284614
rect 354986 248058 355542 248614
rect 354986 212058 355542 212614
rect 354986 176058 355542 176614
rect 354986 140058 355542 140614
rect 354986 104058 355542 104614
rect 354986 68058 355542 68614
rect 354986 32058 355542 32614
rect 336986 -6662 337542 -6106
rect 361826 326898 362382 327454
rect 361826 290898 362382 291454
rect 361826 254898 362382 255454
rect 361826 218898 362382 219454
rect 361826 182898 362382 183454
rect 361826 146898 362382 147454
rect 361826 110898 362382 111454
rect 361826 74898 362382 75454
rect 361826 38898 362382 39454
rect 361826 2898 362382 3454
rect 361826 -902 362382 -346
rect 365546 330618 366102 331174
rect 365546 294618 366102 295174
rect 365546 258618 366102 259174
rect 365546 222618 366102 223174
rect 365546 186618 366102 187174
rect 365546 150618 366102 151174
rect 365546 114618 366102 115174
rect 365546 78618 366102 79174
rect 365546 42618 366102 43174
rect 365546 6618 366102 7174
rect 365546 -2822 366102 -2266
rect 369266 334338 369822 334894
rect 369266 298338 369822 298894
rect 369266 262338 369822 262894
rect 369266 226338 369822 226894
rect 369266 190338 369822 190894
rect 369266 154338 369822 154894
rect 369266 118338 369822 118894
rect 369266 82338 369822 82894
rect 369266 46338 369822 46894
rect 369266 10338 369822 10894
rect 369266 -4742 369822 -4186
rect 372986 302058 373542 302614
rect 372986 266058 373542 266614
rect 372986 230058 373542 230614
rect 372986 194058 373542 194614
rect 372986 158058 373542 158614
rect 372986 122058 373542 122614
rect 372986 86058 373542 86614
rect 372986 50058 373542 50614
rect 372986 14058 373542 14614
rect 354986 -7622 355542 -7066
rect 379826 308898 380382 309454
rect 379826 272898 380382 273454
rect 379826 236898 380382 237454
rect 379826 200898 380382 201454
rect 379826 164898 380382 165454
rect 379826 128898 380382 129454
rect 379826 92898 380382 93454
rect 379826 56898 380382 57454
rect 379826 20898 380382 21454
rect 379826 -1862 380382 -1306
rect 383546 312618 384102 313174
rect 383546 276618 384102 277174
rect 387266 316338 387822 316894
rect 387266 280338 387822 280894
rect 383546 240618 384102 241174
rect 383546 204618 384102 205174
rect 383546 168618 384102 169174
rect 383546 132618 384102 133174
rect 383546 96618 384102 97174
rect 383546 60618 384102 61174
rect 383546 24618 384102 25174
rect 383546 -3782 384102 -3226
rect 392850 435218 393086 435454
rect 392850 434898 393086 435134
rect 392850 399218 393086 399454
rect 392850 398898 393086 399134
rect 392850 363218 393086 363454
rect 392850 362898 393086 363134
rect 390986 320058 391542 320614
rect 390986 284058 391542 284614
rect 387266 244338 387822 244894
rect 390986 248058 391542 248614
rect 387266 208338 387822 208894
rect 387266 172338 387822 172894
rect 387266 136338 387822 136894
rect 387266 100338 387822 100894
rect 387266 64338 387822 64894
rect 387266 28338 387822 28894
rect 387266 -5702 387822 -5146
rect 390986 212058 391542 212614
rect 390986 176058 391542 176614
rect 390986 140058 391542 140614
rect 397826 326898 398382 327454
rect 397826 290898 398382 291454
rect 397826 254898 398382 255454
rect 397826 218898 398382 219454
rect 397826 182898 398382 183454
rect 397826 146898 398382 147454
rect 390986 104058 391542 104614
rect 390986 68058 391542 68614
rect 390986 32058 391542 32614
rect 372986 -6662 373542 -6106
rect 401546 330618 402102 331174
rect 401546 294618 402102 295174
rect 401546 258618 402102 259174
rect 401546 222618 402102 223174
rect 401546 186618 402102 187174
rect 401546 150618 402102 151174
rect 401546 114618 402102 115174
rect 397826 110898 398382 111454
rect 397826 74898 398382 75454
rect 397826 38898 398382 39454
rect 397826 2898 398382 3454
rect 397826 -902 398382 -346
rect 405266 334338 405822 334894
rect 405266 298338 405822 298894
rect 405266 262338 405822 262894
rect 405266 226338 405822 226894
rect 405266 190338 405822 190894
rect 405266 154338 405822 154894
rect 405266 118338 405822 118894
rect 401546 78618 402102 79174
rect 401546 42618 402102 43174
rect 401546 6618 402102 7174
rect 401546 -2822 402102 -2266
rect 405266 82338 405822 82894
rect 408210 453218 408446 453454
rect 408210 452898 408446 453134
rect 408210 417218 408446 417454
rect 408210 416898 408446 417134
rect 408210 381218 408446 381454
rect 408210 380898 408446 381134
rect 408210 345218 408446 345454
rect 408210 344898 408446 345134
rect 408986 302058 409542 302614
rect 408986 266058 409542 266614
rect 408986 230058 409542 230614
rect 408986 194058 409542 194614
rect 408986 158058 409542 158614
rect 408986 122058 409542 122614
rect 408986 86058 409542 86614
rect 405266 46338 405822 46894
rect 405266 10338 405822 10894
rect 405266 -4742 405822 -4186
rect 408986 50058 409542 50614
rect 408986 14058 409542 14614
rect 390986 -7622 391542 -7066
rect 415826 452898 416382 453454
rect 415826 416898 416382 417454
rect 415826 380898 416382 381454
rect 415826 344898 416382 345454
rect 415826 308898 416382 309454
rect 415826 272898 416382 273454
rect 415826 236898 416382 237454
rect 415826 200898 416382 201454
rect 415826 164898 416382 165454
rect 415826 128898 416382 129454
rect 415826 92898 416382 93454
rect 415826 56898 416382 57454
rect 415826 20898 416382 21454
rect 415826 -1862 416382 -1306
rect 419546 672618 420102 673174
rect 419546 636618 420102 637174
rect 419546 600618 420102 601174
rect 419546 564618 420102 565174
rect 419546 528618 420102 529174
rect 419546 492618 420102 493174
rect 419546 456618 420102 457174
rect 419546 420618 420102 421174
rect 419546 384618 420102 385174
rect 419546 348618 420102 349174
rect 419546 312618 420102 313174
rect 419546 276618 420102 277174
rect 419546 240618 420102 241174
rect 419546 204618 420102 205174
rect 419546 168618 420102 169174
rect 419546 132618 420102 133174
rect 419546 96618 420102 97174
rect 419546 60618 420102 61174
rect 419546 24618 420102 25174
rect 419546 -3782 420102 -3226
rect 423266 676338 423822 676894
rect 423266 640338 423822 640894
rect 423266 604338 423822 604894
rect 423266 568338 423822 568894
rect 423266 532338 423822 532894
rect 423266 496338 423822 496894
rect 423266 460338 423822 460894
rect 423266 424338 423822 424894
rect 423266 388338 423822 388894
rect 423266 352338 423822 352894
rect 423266 316338 423822 316894
rect 423266 280338 423822 280894
rect 423266 244338 423822 244894
rect 423266 208338 423822 208894
rect 423266 172338 423822 172894
rect 423266 136338 423822 136894
rect 423266 100338 423822 100894
rect 423266 64338 423822 64894
rect 423266 28338 423822 28894
rect 423266 -5702 423822 -5146
rect 444986 710042 445542 710598
rect 441266 708122 441822 708678
rect 437546 706202 438102 706758
rect 426986 680058 427542 680614
rect 426986 644058 427542 644614
rect 426986 608058 427542 608614
rect 426986 572058 427542 572614
rect 426986 536058 427542 536614
rect 426986 500058 427542 500614
rect 426986 464058 427542 464614
rect 426986 428058 427542 428614
rect 426986 392058 427542 392614
rect 426986 356058 427542 356614
rect 426986 320058 427542 320614
rect 426986 284058 427542 284614
rect 426986 248058 427542 248614
rect 426986 212058 427542 212614
rect 426986 176058 427542 176614
rect 426986 140058 427542 140614
rect 426986 104058 427542 104614
rect 426986 68058 427542 68614
rect 426986 32058 427542 32614
rect 408986 -6662 409542 -6106
rect 433826 704282 434382 704838
rect 433826 686898 434382 687454
rect 433826 650898 434382 651454
rect 433826 614898 434382 615454
rect 433826 578898 434382 579454
rect 433826 542898 434382 543454
rect 433826 506898 434382 507454
rect 433826 470898 434382 471454
rect 433826 434898 434382 435454
rect 433826 398898 434382 399454
rect 433826 362898 434382 363454
rect 433826 326898 434382 327454
rect 433826 290898 434382 291454
rect 433826 254898 434382 255454
rect 433826 218898 434382 219454
rect 433826 182898 434382 183454
rect 433826 146898 434382 147454
rect 433826 110898 434382 111454
rect 433826 74898 434382 75454
rect 433826 38898 434382 39454
rect 433826 2898 434382 3454
rect 433826 -902 434382 -346
rect 437546 690618 438102 691174
rect 437546 654618 438102 655174
rect 437546 618618 438102 619174
rect 437546 582618 438102 583174
rect 437546 546618 438102 547174
rect 437546 510618 438102 511174
rect 437546 474618 438102 475174
rect 437546 438618 438102 439174
rect 437546 402618 438102 403174
rect 437546 366618 438102 367174
rect 437546 330618 438102 331174
rect 437546 294618 438102 295174
rect 437546 258618 438102 259174
rect 437546 222618 438102 223174
rect 437546 186618 438102 187174
rect 437546 150618 438102 151174
rect 437546 114618 438102 115174
rect 437546 78618 438102 79174
rect 437546 42618 438102 43174
rect 437546 6618 438102 7174
rect 437546 -2822 438102 -2266
rect 441266 694338 441822 694894
rect 441266 658338 441822 658894
rect 441266 622338 441822 622894
rect 441266 586338 441822 586894
rect 441266 550338 441822 550894
rect 441266 514338 441822 514894
rect 441266 478338 441822 478894
rect 441266 442338 441822 442894
rect 441266 406338 441822 406894
rect 441266 370338 441822 370894
rect 441266 334338 441822 334894
rect 441266 298338 441822 298894
rect 441266 262338 441822 262894
rect 441266 226338 441822 226894
rect 441266 190338 441822 190894
rect 441266 154338 441822 154894
rect 441266 118338 441822 118894
rect 441266 82338 441822 82894
rect 441266 46338 441822 46894
rect 441266 10338 441822 10894
rect 441266 -4742 441822 -4186
rect 462986 711002 463542 711558
rect 459266 709082 459822 709638
rect 455546 707162 456102 707718
rect 444986 698058 445542 698614
rect 444986 662058 445542 662614
rect 444986 626058 445542 626614
rect 444986 590058 445542 590614
rect 444986 554058 445542 554614
rect 444986 518058 445542 518614
rect 444986 482058 445542 482614
rect 444986 446058 445542 446614
rect 444986 410058 445542 410614
rect 444986 374058 445542 374614
rect 444986 338058 445542 338614
rect 444986 302058 445542 302614
rect 444986 266058 445542 266614
rect 444986 230058 445542 230614
rect 444986 194058 445542 194614
rect 444986 158058 445542 158614
rect 444986 122058 445542 122614
rect 444986 86058 445542 86614
rect 444986 50058 445542 50614
rect 444986 14058 445542 14614
rect 426986 -7622 427542 -7066
rect 451826 705242 452382 705798
rect 451826 668898 452382 669454
rect 451826 632898 452382 633454
rect 451826 596898 452382 597454
rect 451826 560898 452382 561454
rect 451826 524898 452382 525454
rect 451826 488898 452382 489454
rect 451826 452898 452382 453454
rect 451826 416898 452382 417454
rect 451826 380898 452382 381454
rect 451826 344898 452382 345454
rect 451826 308898 452382 309454
rect 451826 272898 452382 273454
rect 451826 236898 452382 237454
rect 451826 200898 452382 201454
rect 451826 164898 452382 165454
rect 451826 128898 452382 129454
rect 451826 92898 452382 93454
rect 451826 56898 452382 57454
rect 451826 20898 452382 21454
rect 451826 -1862 452382 -1306
rect 455546 672618 456102 673174
rect 455546 636618 456102 637174
rect 455546 600618 456102 601174
rect 455546 564618 456102 565174
rect 455546 528618 456102 529174
rect 455546 492618 456102 493174
rect 455546 456618 456102 457174
rect 455546 420618 456102 421174
rect 455546 384618 456102 385174
rect 455546 348618 456102 349174
rect 455546 312618 456102 313174
rect 455546 276618 456102 277174
rect 455546 240618 456102 241174
rect 455546 204618 456102 205174
rect 455546 168618 456102 169174
rect 455546 132618 456102 133174
rect 455546 96618 456102 97174
rect 455546 60618 456102 61174
rect 455546 24618 456102 25174
rect 455546 -3782 456102 -3226
rect 459266 676338 459822 676894
rect 459266 640338 459822 640894
rect 459266 604338 459822 604894
rect 459266 568338 459822 568894
rect 459266 532338 459822 532894
rect 459266 496338 459822 496894
rect 459266 460338 459822 460894
rect 459266 424338 459822 424894
rect 459266 388338 459822 388894
rect 459266 352338 459822 352894
rect 459266 316338 459822 316894
rect 459266 280338 459822 280894
rect 459266 244338 459822 244894
rect 459266 208338 459822 208894
rect 459266 172338 459822 172894
rect 459266 136338 459822 136894
rect 459266 100338 459822 100894
rect 459266 64338 459822 64894
rect 459266 28338 459822 28894
rect 459266 -5702 459822 -5146
rect 480986 710042 481542 710598
rect 477266 708122 477822 708678
rect 473546 706202 474102 706758
rect 462986 680058 463542 680614
rect 462986 644058 463542 644614
rect 462986 608058 463542 608614
rect 462986 572058 463542 572614
rect 462986 536058 463542 536614
rect 462986 500058 463542 500614
rect 462986 464058 463542 464614
rect 462986 428058 463542 428614
rect 462986 392058 463542 392614
rect 462986 356058 463542 356614
rect 462986 320058 463542 320614
rect 462986 284058 463542 284614
rect 462986 248058 463542 248614
rect 462986 212058 463542 212614
rect 462986 176058 463542 176614
rect 462986 140058 463542 140614
rect 462986 104058 463542 104614
rect 462986 68058 463542 68614
rect 462986 32058 463542 32614
rect 444986 -6662 445542 -6106
rect 469826 704282 470382 704838
rect 469826 686898 470382 687454
rect 469826 650898 470382 651454
rect 469826 614898 470382 615454
rect 469826 578898 470382 579454
rect 469826 542898 470382 543454
rect 469826 506898 470382 507454
rect 469826 470898 470382 471454
rect 469826 434898 470382 435454
rect 469826 398898 470382 399454
rect 469826 362898 470382 363454
rect 469826 326898 470382 327454
rect 469826 290898 470382 291454
rect 469826 254898 470382 255454
rect 469826 218898 470382 219454
rect 469826 182898 470382 183454
rect 469826 146898 470382 147454
rect 469826 110898 470382 111454
rect 469826 74898 470382 75454
rect 469826 38898 470382 39454
rect 469826 2898 470382 3454
rect 469826 -902 470382 -346
rect 473546 690618 474102 691174
rect 473546 654618 474102 655174
rect 473546 618618 474102 619174
rect 473546 582618 474102 583174
rect 473546 546618 474102 547174
rect 473546 510618 474102 511174
rect 473546 474618 474102 475174
rect 473546 438618 474102 439174
rect 473546 402618 474102 403174
rect 473546 366618 474102 367174
rect 473546 330618 474102 331174
rect 473546 294618 474102 295174
rect 473546 258618 474102 259174
rect 473546 222618 474102 223174
rect 473546 186618 474102 187174
rect 473546 150618 474102 151174
rect 473546 114618 474102 115174
rect 473546 78618 474102 79174
rect 473546 42618 474102 43174
rect 473546 6618 474102 7174
rect 473546 -2822 474102 -2266
rect 477266 694338 477822 694894
rect 477266 658338 477822 658894
rect 477266 622338 477822 622894
rect 477266 586338 477822 586894
rect 477266 550338 477822 550894
rect 477266 514338 477822 514894
rect 477266 478338 477822 478894
rect 477266 442338 477822 442894
rect 477266 406338 477822 406894
rect 477266 370338 477822 370894
rect 477266 334338 477822 334894
rect 477266 298338 477822 298894
rect 477266 262338 477822 262894
rect 477266 226338 477822 226894
rect 477266 190338 477822 190894
rect 477266 154338 477822 154894
rect 477266 118338 477822 118894
rect 477266 82338 477822 82894
rect 477266 46338 477822 46894
rect 477266 10338 477822 10894
rect 477266 -4742 477822 -4186
rect 498986 711002 499542 711558
rect 495266 709082 495822 709638
rect 491546 707162 492102 707718
rect 480986 698058 481542 698614
rect 480986 662058 481542 662614
rect 480986 626058 481542 626614
rect 480986 590058 481542 590614
rect 480986 554058 481542 554614
rect 480986 518058 481542 518614
rect 480986 482058 481542 482614
rect 480986 446058 481542 446614
rect 480986 410058 481542 410614
rect 480986 374058 481542 374614
rect 480986 338058 481542 338614
rect 480986 302058 481542 302614
rect 480986 266058 481542 266614
rect 480986 230058 481542 230614
rect 480986 194058 481542 194614
rect 480986 158058 481542 158614
rect 480986 122058 481542 122614
rect 480986 86058 481542 86614
rect 480986 50058 481542 50614
rect 480986 14058 481542 14614
rect 462986 -7622 463542 -7066
rect 487826 705242 488382 705798
rect 487826 668898 488382 669454
rect 487826 632898 488382 633454
rect 487826 596898 488382 597454
rect 487826 560898 488382 561454
rect 487826 524898 488382 525454
rect 487826 488898 488382 489454
rect 487826 452898 488382 453454
rect 487826 416898 488382 417454
rect 487826 380898 488382 381454
rect 487826 344898 488382 345454
rect 487826 308898 488382 309454
rect 487826 272898 488382 273454
rect 487826 236898 488382 237454
rect 487826 200898 488382 201454
rect 487826 164898 488382 165454
rect 487826 128898 488382 129454
rect 487826 92898 488382 93454
rect 487826 56898 488382 57454
rect 487826 20898 488382 21454
rect 487826 -1862 488382 -1306
rect 491546 672618 492102 673174
rect 491546 636618 492102 637174
rect 491546 600618 492102 601174
rect 491546 564618 492102 565174
rect 491546 528618 492102 529174
rect 491546 492618 492102 493174
rect 491546 456618 492102 457174
rect 491546 420618 492102 421174
rect 491546 384618 492102 385174
rect 491546 348618 492102 349174
rect 491546 312618 492102 313174
rect 491546 276618 492102 277174
rect 491546 240618 492102 241174
rect 491546 204618 492102 205174
rect 491546 168618 492102 169174
rect 491546 132618 492102 133174
rect 491546 96618 492102 97174
rect 491546 60618 492102 61174
rect 491546 24618 492102 25174
rect 491546 -3782 492102 -3226
rect 495266 676338 495822 676894
rect 495266 640338 495822 640894
rect 495266 604338 495822 604894
rect 495266 568338 495822 568894
rect 495266 532338 495822 532894
rect 495266 496338 495822 496894
rect 495266 460338 495822 460894
rect 495266 424338 495822 424894
rect 495266 388338 495822 388894
rect 495266 352338 495822 352894
rect 495266 316338 495822 316894
rect 495266 280338 495822 280894
rect 495266 244338 495822 244894
rect 495266 208338 495822 208894
rect 495266 172338 495822 172894
rect 495266 136338 495822 136894
rect 495266 100338 495822 100894
rect 495266 64338 495822 64894
rect 495266 28338 495822 28894
rect 495266 -5702 495822 -5146
rect 516986 710042 517542 710598
rect 513266 708122 513822 708678
rect 509546 706202 510102 706758
rect 498986 680058 499542 680614
rect 498986 644058 499542 644614
rect 498986 608058 499542 608614
rect 498986 572058 499542 572614
rect 498986 536058 499542 536614
rect 498986 500058 499542 500614
rect 498986 464058 499542 464614
rect 498986 428058 499542 428614
rect 498986 392058 499542 392614
rect 498986 356058 499542 356614
rect 498986 320058 499542 320614
rect 498986 284058 499542 284614
rect 498986 248058 499542 248614
rect 498986 212058 499542 212614
rect 498986 176058 499542 176614
rect 498986 140058 499542 140614
rect 498986 104058 499542 104614
rect 498986 68058 499542 68614
rect 498986 32058 499542 32614
rect 480986 -6662 481542 -6106
rect 505826 704282 506382 704838
rect 505826 686898 506382 687454
rect 505826 650898 506382 651454
rect 505826 614898 506382 615454
rect 505826 578898 506382 579454
rect 505826 542898 506382 543454
rect 505826 506898 506382 507454
rect 505826 470898 506382 471454
rect 505826 434898 506382 435454
rect 505826 398898 506382 399454
rect 505826 362898 506382 363454
rect 505826 326898 506382 327454
rect 505826 290898 506382 291454
rect 505826 254898 506382 255454
rect 505826 218898 506382 219454
rect 505826 182898 506382 183454
rect 505826 146898 506382 147454
rect 505826 110898 506382 111454
rect 505826 74898 506382 75454
rect 505826 38898 506382 39454
rect 505826 2898 506382 3454
rect 505826 -902 506382 -346
rect 509546 690618 510102 691174
rect 509546 654618 510102 655174
rect 509546 618618 510102 619174
rect 509546 582618 510102 583174
rect 509546 546618 510102 547174
rect 509546 510618 510102 511174
rect 509546 474618 510102 475174
rect 509546 438618 510102 439174
rect 509546 402618 510102 403174
rect 509546 366618 510102 367174
rect 509546 330618 510102 331174
rect 509546 294618 510102 295174
rect 509546 258618 510102 259174
rect 509546 222618 510102 223174
rect 509546 186618 510102 187174
rect 509546 150618 510102 151174
rect 509546 114618 510102 115174
rect 509546 78618 510102 79174
rect 509546 42618 510102 43174
rect 509546 6618 510102 7174
rect 509546 -2822 510102 -2266
rect 513266 694338 513822 694894
rect 513266 658338 513822 658894
rect 513266 622338 513822 622894
rect 513266 586338 513822 586894
rect 513266 550338 513822 550894
rect 513266 514338 513822 514894
rect 513266 478338 513822 478894
rect 513266 442338 513822 442894
rect 513266 406338 513822 406894
rect 513266 370338 513822 370894
rect 513266 334338 513822 334894
rect 513266 298338 513822 298894
rect 513266 262338 513822 262894
rect 513266 226338 513822 226894
rect 513266 190338 513822 190894
rect 513266 154338 513822 154894
rect 513266 118338 513822 118894
rect 513266 82338 513822 82894
rect 513266 46338 513822 46894
rect 513266 10338 513822 10894
rect 513266 -4742 513822 -4186
rect 534986 711002 535542 711558
rect 531266 709082 531822 709638
rect 527546 707162 528102 707718
rect 516986 698058 517542 698614
rect 516986 662058 517542 662614
rect 516986 626058 517542 626614
rect 516986 590058 517542 590614
rect 516986 554058 517542 554614
rect 516986 518058 517542 518614
rect 516986 482058 517542 482614
rect 516986 446058 517542 446614
rect 516986 410058 517542 410614
rect 516986 374058 517542 374614
rect 516986 338058 517542 338614
rect 516986 302058 517542 302614
rect 516986 266058 517542 266614
rect 516986 230058 517542 230614
rect 516986 194058 517542 194614
rect 516986 158058 517542 158614
rect 516986 122058 517542 122614
rect 516986 86058 517542 86614
rect 516986 50058 517542 50614
rect 516986 14058 517542 14614
rect 498986 -7622 499542 -7066
rect 523826 705242 524382 705798
rect 523826 668898 524382 669454
rect 523826 632898 524382 633454
rect 523826 596898 524382 597454
rect 523826 560898 524382 561454
rect 523826 524898 524382 525454
rect 523826 488898 524382 489454
rect 523826 452898 524382 453454
rect 523826 416898 524382 417454
rect 523826 380898 524382 381454
rect 523826 344898 524382 345454
rect 523826 308898 524382 309454
rect 523826 272898 524382 273454
rect 523826 236898 524382 237454
rect 523826 200898 524382 201454
rect 523826 164898 524382 165454
rect 523826 128898 524382 129454
rect 523826 92898 524382 93454
rect 523826 56898 524382 57454
rect 523826 20898 524382 21454
rect 523826 -1862 524382 -1306
rect 527546 672618 528102 673174
rect 527546 636618 528102 637174
rect 527546 600618 528102 601174
rect 527546 564618 528102 565174
rect 527546 528618 528102 529174
rect 527546 492618 528102 493174
rect 527546 456618 528102 457174
rect 527546 420618 528102 421174
rect 527546 384618 528102 385174
rect 527546 348618 528102 349174
rect 527546 312618 528102 313174
rect 527546 276618 528102 277174
rect 527546 240618 528102 241174
rect 527546 204618 528102 205174
rect 527546 168618 528102 169174
rect 527546 132618 528102 133174
rect 527546 96618 528102 97174
rect 527546 60618 528102 61174
rect 527546 24618 528102 25174
rect 527546 -3782 528102 -3226
rect 531266 676338 531822 676894
rect 531266 640338 531822 640894
rect 531266 604338 531822 604894
rect 531266 568338 531822 568894
rect 531266 532338 531822 532894
rect 531266 496338 531822 496894
rect 531266 460338 531822 460894
rect 531266 424338 531822 424894
rect 531266 388338 531822 388894
rect 531266 352338 531822 352894
rect 531266 316338 531822 316894
rect 531266 280338 531822 280894
rect 531266 244338 531822 244894
rect 531266 208338 531822 208894
rect 531266 172338 531822 172894
rect 531266 136338 531822 136894
rect 531266 100338 531822 100894
rect 531266 64338 531822 64894
rect 531266 28338 531822 28894
rect 531266 -5702 531822 -5146
rect 552986 710042 553542 710598
rect 549266 708122 549822 708678
rect 545546 706202 546102 706758
rect 534986 680058 535542 680614
rect 534986 644058 535542 644614
rect 534986 608058 535542 608614
rect 534986 572058 535542 572614
rect 534986 536058 535542 536614
rect 534986 500058 535542 500614
rect 534986 464058 535542 464614
rect 534986 428058 535542 428614
rect 534986 392058 535542 392614
rect 534986 356058 535542 356614
rect 534986 320058 535542 320614
rect 534986 284058 535542 284614
rect 534986 248058 535542 248614
rect 534986 212058 535542 212614
rect 534986 176058 535542 176614
rect 534986 140058 535542 140614
rect 534986 104058 535542 104614
rect 534986 68058 535542 68614
rect 534986 32058 535542 32614
rect 516986 -6662 517542 -6106
rect 541826 704282 542382 704838
rect 541826 686898 542382 687454
rect 541826 650898 542382 651454
rect 541826 614898 542382 615454
rect 541826 578898 542382 579454
rect 541826 542898 542382 543454
rect 541826 506898 542382 507454
rect 541826 470898 542382 471454
rect 541826 434898 542382 435454
rect 541826 398898 542382 399454
rect 541826 362898 542382 363454
rect 541826 326898 542382 327454
rect 541826 290898 542382 291454
rect 541826 254898 542382 255454
rect 541826 218898 542382 219454
rect 541826 182898 542382 183454
rect 541826 146898 542382 147454
rect 541826 110898 542382 111454
rect 541826 74898 542382 75454
rect 541826 38898 542382 39454
rect 541826 2898 542382 3454
rect 541826 -902 542382 -346
rect 545546 690618 546102 691174
rect 545546 654618 546102 655174
rect 545546 618618 546102 619174
rect 545546 582618 546102 583174
rect 545546 546618 546102 547174
rect 545546 510618 546102 511174
rect 545546 474618 546102 475174
rect 545546 438618 546102 439174
rect 545546 402618 546102 403174
rect 545546 366618 546102 367174
rect 545546 330618 546102 331174
rect 545546 294618 546102 295174
rect 545546 258618 546102 259174
rect 545546 222618 546102 223174
rect 545546 186618 546102 187174
rect 545546 150618 546102 151174
rect 545546 114618 546102 115174
rect 545546 78618 546102 79174
rect 545546 42618 546102 43174
rect 545546 6618 546102 7174
rect 545546 -2822 546102 -2266
rect 549266 694338 549822 694894
rect 549266 658338 549822 658894
rect 549266 622338 549822 622894
rect 549266 586338 549822 586894
rect 549266 550338 549822 550894
rect 549266 514338 549822 514894
rect 549266 478338 549822 478894
rect 549266 442338 549822 442894
rect 549266 406338 549822 406894
rect 549266 370338 549822 370894
rect 549266 334338 549822 334894
rect 549266 298338 549822 298894
rect 549266 262338 549822 262894
rect 549266 226338 549822 226894
rect 549266 190338 549822 190894
rect 549266 154338 549822 154894
rect 549266 118338 549822 118894
rect 549266 82338 549822 82894
rect 549266 46338 549822 46894
rect 549266 10338 549822 10894
rect 549266 -4742 549822 -4186
rect 570986 711002 571542 711558
rect 567266 709082 567822 709638
rect 563546 707162 564102 707718
rect 552986 698058 553542 698614
rect 552986 662058 553542 662614
rect 552986 626058 553542 626614
rect 552986 590058 553542 590614
rect 552986 554058 553542 554614
rect 552986 518058 553542 518614
rect 552986 482058 553542 482614
rect 552986 446058 553542 446614
rect 552986 410058 553542 410614
rect 552986 374058 553542 374614
rect 552986 338058 553542 338614
rect 552986 302058 553542 302614
rect 552986 266058 553542 266614
rect 552986 230058 553542 230614
rect 552986 194058 553542 194614
rect 552986 158058 553542 158614
rect 552986 122058 553542 122614
rect 552986 86058 553542 86614
rect 552986 50058 553542 50614
rect 552986 14058 553542 14614
rect 534986 -7622 535542 -7066
rect 559826 705242 560382 705798
rect 559826 668898 560382 669454
rect 559826 632898 560382 633454
rect 559826 596898 560382 597454
rect 559826 560898 560382 561454
rect 559826 524898 560382 525454
rect 559826 488898 560382 489454
rect 559826 452898 560382 453454
rect 559826 416898 560382 417454
rect 559826 380898 560382 381454
rect 559826 344898 560382 345454
rect 559826 308898 560382 309454
rect 559826 272898 560382 273454
rect 559826 236898 560382 237454
rect 559826 200898 560382 201454
rect 559826 164898 560382 165454
rect 559826 128898 560382 129454
rect 559826 92898 560382 93454
rect 559826 56898 560382 57454
rect 559826 20898 560382 21454
rect 559826 -1862 560382 -1306
rect 563546 672618 564102 673174
rect 563546 636618 564102 637174
rect 563546 600618 564102 601174
rect 563546 564618 564102 565174
rect 563546 528618 564102 529174
rect 563546 492618 564102 493174
rect 563546 456618 564102 457174
rect 563546 420618 564102 421174
rect 563546 384618 564102 385174
rect 563546 348618 564102 349174
rect 563546 312618 564102 313174
rect 563546 276618 564102 277174
rect 563546 240618 564102 241174
rect 563546 204618 564102 205174
rect 563546 168618 564102 169174
rect 563546 132618 564102 133174
rect 563546 96618 564102 97174
rect 563546 60618 564102 61174
rect 563546 24618 564102 25174
rect 563546 -3782 564102 -3226
rect 567266 676338 567822 676894
rect 567266 640338 567822 640894
rect 567266 604338 567822 604894
rect 567266 568338 567822 568894
rect 567266 532338 567822 532894
rect 567266 496338 567822 496894
rect 567266 460338 567822 460894
rect 567266 424338 567822 424894
rect 567266 388338 567822 388894
rect 567266 352338 567822 352894
rect 567266 316338 567822 316894
rect 567266 280338 567822 280894
rect 567266 244338 567822 244894
rect 567266 208338 567822 208894
rect 567266 172338 567822 172894
rect 567266 136338 567822 136894
rect 567266 100338 567822 100894
rect 567266 64338 567822 64894
rect 567266 28338 567822 28894
rect 567266 -5702 567822 -5146
rect 592062 711002 592618 711558
rect 591102 710042 591658 710598
rect 590142 709082 590698 709638
rect 589182 708122 589738 708678
rect 588222 707162 588778 707718
rect 581546 706202 582102 706758
rect 570986 680058 571542 680614
rect 570986 644058 571542 644614
rect 570986 608058 571542 608614
rect 570986 572058 571542 572614
rect 570986 536058 571542 536614
rect 570986 500058 571542 500614
rect 570986 464058 571542 464614
rect 570986 428058 571542 428614
rect 570986 392058 571542 392614
rect 570986 356058 571542 356614
rect 570986 320058 571542 320614
rect 570986 284058 571542 284614
rect 570986 248058 571542 248614
rect 570986 212058 571542 212614
rect 570986 176058 571542 176614
rect 570986 140058 571542 140614
rect 570986 104058 571542 104614
rect 570986 68058 571542 68614
rect 570986 32058 571542 32614
rect 552986 -6662 553542 -6106
rect 577826 704282 578382 704838
rect 577826 686898 578382 687454
rect 577826 650898 578382 651454
rect 577826 614898 578382 615454
rect 577826 578898 578382 579454
rect 577826 542898 578382 543454
rect 577826 506898 578382 507454
rect 577826 470898 578382 471454
rect 577826 434898 578382 435454
rect 577826 398898 578382 399454
rect 577826 362898 578382 363454
rect 577826 326898 578382 327454
rect 577826 290898 578382 291454
rect 577826 254898 578382 255454
rect 577826 218898 578382 219454
rect 577826 182898 578382 183454
rect 577826 146898 578382 147454
rect 577826 110898 578382 111454
rect 577826 74898 578382 75454
rect 577826 38898 578382 39454
rect 577826 2898 578382 3454
rect 577826 -902 578382 -346
rect 587262 706202 587818 706758
rect 586302 705242 586858 705798
rect 581546 690618 582102 691174
rect 581546 654618 582102 655174
rect 581546 618618 582102 619174
rect 581546 582618 582102 583174
rect 581546 546618 582102 547174
rect 581546 510618 582102 511174
rect 581546 474618 582102 475174
rect 581546 438618 582102 439174
rect 581546 402618 582102 403174
rect 581546 366618 582102 367174
rect 581546 330618 582102 331174
rect 581546 294618 582102 295174
rect 581546 258618 582102 259174
rect 581546 222618 582102 223174
rect 581546 186618 582102 187174
rect 581546 150618 582102 151174
rect 581546 114618 582102 115174
rect 581546 78618 582102 79174
rect 581546 42618 582102 43174
rect 581546 6618 582102 7174
rect 585342 704282 585898 704838
rect 585342 686898 585898 687454
rect 585342 650898 585898 651454
rect 585342 614898 585898 615454
rect 585342 578898 585898 579454
rect 585342 542898 585898 543454
rect 585342 506898 585898 507454
rect 585342 470898 585898 471454
rect 585342 434898 585898 435454
rect 585342 398898 585898 399454
rect 585342 362898 585898 363454
rect 585342 326898 585898 327454
rect 585342 290898 585898 291454
rect 585342 254898 585898 255454
rect 585342 218898 585898 219454
rect 585342 182898 585898 183454
rect 585342 146898 585898 147454
rect 585342 110898 585898 111454
rect 585342 74898 585898 75454
rect 585342 38898 585898 39454
rect 585342 2898 585898 3454
rect 585342 -902 585898 -346
rect 586302 668898 586858 669454
rect 586302 632898 586858 633454
rect 586302 596898 586858 597454
rect 586302 560898 586858 561454
rect 586302 524898 586858 525454
rect 586302 488898 586858 489454
rect 586302 452898 586858 453454
rect 586302 416898 586858 417454
rect 586302 380898 586858 381454
rect 586302 344898 586858 345454
rect 586302 308898 586858 309454
rect 586302 272898 586858 273454
rect 586302 236898 586858 237454
rect 586302 200898 586858 201454
rect 586302 164898 586858 165454
rect 586302 128898 586858 129454
rect 586302 92898 586858 93454
rect 586302 56898 586858 57454
rect 586302 20898 586858 21454
rect 586302 -1862 586858 -1306
rect 587262 690618 587818 691174
rect 587262 654618 587818 655174
rect 587262 618618 587818 619174
rect 587262 582618 587818 583174
rect 587262 546618 587818 547174
rect 587262 510618 587818 511174
rect 587262 474618 587818 475174
rect 587262 438618 587818 439174
rect 587262 402618 587818 403174
rect 587262 366618 587818 367174
rect 587262 330618 587818 331174
rect 587262 294618 587818 295174
rect 587262 258618 587818 259174
rect 587262 222618 587818 223174
rect 587262 186618 587818 187174
rect 587262 150618 587818 151174
rect 587262 114618 587818 115174
rect 587262 78618 587818 79174
rect 587262 42618 587818 43174
rect 587262 6618 587818 7174
rect 581546 -2822 582102 -2266
rect 587262 -2822 587818 -2266
rect 588222 672618 588778 673174
rect 588222 636618 588778 637174
rect 588222 600618 588778 601174
rect 588222 564618 588778 565174
rect 588222 528618 588778 529174
rect 588222 492618 588778 493174
rect 588222 456618 588778 457174
rect 588222 420618 588778 421174
rect 588222 384618 588778 385174
rect 588222 348618 588778 349174
rect 588222 312618 588778 313174
rect 588222 276618 588778 277174
rect 588222 240618 588778 241174
rect 588222 204618 588778 205174
rect 588222 168618 588778 169174
rect 588222 132618 588778 133174
rect 588222 96618 588778 97174
rect 588222 60618 588778 61174
rect 588222 24618 588778 25174
rect 588222 -3782 588778 -3226
rect 589182 694338 589738 694894
rect 589182 658338 589738 658894
rect 589182 622338 589738 622894
rect 589182 586338 589738 586894
rect 589182 550338 589738 550894
rect 589182 514338 589738 514894
rect 589182 478338 589738 478894
rect 589182 442338 589738 442894
rect 589182 406338 589738 406894
rect 589182 370338 589738 370894
rect 589182 334338 589738 334894
rect 589182 298338 589738 298894
rect 589182 262338 589738 262894
rect 589182 226338 589738 226894
rect 589182 190338 589738 190894
rect 589182 154338 589738 154894
rect 589182 118338 589738 118894
rect 589182 82338 589738 82894
rect 589182 46338 589738 46894
rect 589182 10338 589738 10894
rect 589182 -4742 589738 -4186
rect 590142 676338 590698 676894
rect 590142 640338 590698 640894
rect 590142 604338 590698 604894
rect 590142 568338 590698 568894
rect 590142 532338 590698 532894
rect 590142 496338 590698 496894
rect 590142 460338 590698 460894
rect 590142 424338 590698 424894
rect 590142 388338 590698 388894
rect 590142 352338 590698 352894
rect 590142 316338 590698 316894
rect 590142 280338 590698 280894
rect 590142 244338 590698 244894
rect 590142 208338 590698 208894
rect 590142 172338 590698 172894
rect 590142 136338 590698 136894
rect 590142 100338 590698 100894
rect 590142 64338 590698 64894
rect 590142 28338 590698 28894
rect 590142 -5702 590698 -5146
rect 591102 698058 591658 698614
rect 591102 662058 591658 662614
rect 591102 626058 591658 626614
rect 591102 590058 591658 590614
rect 591102 554058 591658 554614
rect 591102 518058 591658 518614
rect 591102 482058 591658 482614
rect 591102 446058 591658 446614
rect 591102 410058 591658 410614
rect 591102 374058 591658 374614
rect 591102 338058 591658 338614
rect 591102 302058 591658 302614
rect 591102 266058 591658 266614
rect 591102 230058 591658 230614
rect 591102 194058 591658 194614
rect 591102 158058 591658 158614
rect 591102 122058 591658 122614
rect 591102 86058 591658 86614
rect 591102 50058 591658 50614
rect 591102 14058 591658 14614
rect 591102 -6662 591658 -6106
rect 592062 680058 592618 680614
rect 592062 644058 592618 644614
rect 592062 608058 592618 608614
rect 592062 572058 592618 572614
rect 592062 536058 592618 536614
rect 592062 500058 592618 500614
rect 592062 464058 592618 464614
rect 592062 428058 592618 428614
rect 592062 392058 592618 392614
rect 592062 356058 592618 356614
rect 592062 320058 592618 320614
rect 592062 284058 592618 284614
rect 592062 248058 592618 248614
rect 592062 212058 592618 212614
rect 592062 176058 592618 176614
rect 592062 140058 592618 140614
rect 592062 104058 592618 104614
rect 592062 68058 592618 68614
rect 592062 32058 592618 32614
rect 570986 -7622 571542 -7066
rect 592062 -7622 592618 -7066
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711002 -8694 711558
rect -8138 711002 30986 711558
rect 31542 711002 66986 711558
rect 67542 711002 102986 711558
rect 103542 711002 138986 711558
rect 139542 711002 174986 711558
rect 175542 711002 210986 711558
rect 211542 711002 246986 711558
rect 247542 711002 282986 711558
rect 283542 711002 318986 711558
rect 319542 711002 354986 711558
rect 355542 711002 390986 711558
rect 391542 711002 426986 711558
rect 427542 711002 462986 711558
rect 463542 711002 498986 711558
rect 499542 711002 534986 711558
rect 535542 711002 570986 711558
rect 571542 711002 592062 711558
rect 592618 711002 592650 711558
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710042 -7734 710598
rect -7178 710042 12986 710598
rect 13542 710042 48986 710598
rect 49542 710042 84986 710598
rect 85542 710042 120986 710598
rect 121542 710042 156986 710598
rect 157542 710042 192986 710598
rect 193542 710042 228986 710598
rect 229542 710042 264986 710598
rect 265542 710042 300986 710598
rect 301542 710042 336986 710598
rect 337542 710042 372986 710598
rect 373542 710042 408986 710598
rect 409542 710042 444986 710598
rect 445542 710042 480986 710598
rect 481542 710042 516986 710598
rect 517542 710042 552986 710598
rect 553542 710042 591102 710598
rect 591658 710042 591690 710598
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709082 -6774 709638
rect -6218 709082 27266 709638
rect 27822 709082 63266 709638
rect 63822 709082 99266 709638
rect 99822 709082 135266 709638
rect 135822 709082 171266 709638
rect 171822 709082 207266 709638
rect 207822 709082 243266 709638
rect 243822 709082 279266 709638
rect 279822 709082 315266 709638
rect 315822 709082 351266 709638
rect 351822 709082 387266 709638
rect 387822 709082 423266 709638
rect 423822 709082 459266 709638
rect 459822 709082 495266 709638
rect 495822 709082 531266 709638
rect 531822 709082 567266 709638
rect 567822 709082 590142 709638
rect 590698 709082 590730 709638
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708122 -5814 708678
rect -5258 708122 9266 708678
rect 9822 708122 45266 708678
rect 45822 708122 81266 708678
rect 81822 708122 117266 708678
rect 117822 708122 153266 708678
rect 153822 708122 189266 708678
rect 189822 708122 225266 708678
rect 225822 708122 261266 708678
rect 261822 708122 297266 708678
rect 297822 708122 333266 708678
rect 333822 708122 369266 708678
rect 369822 708122 405266 708678
rect 405822 708122 441266 708678
rect 441822 708122 477266 708678
rect 477822 708122 513266 708678
rect 513822 708122 549266 708678
rect 549822 708122 589182 708678
rect 589738 708122 589770 708678
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707162 -4854 707718
rect -4298 707162 23546 707718
rect 24102 707162 59546 707718
rect 60102 707162 95546 707718
rect 96102 707162 131546 707718
rect 132102 707162 167546 707718
rect 168102 707162 203546 707718
rect 204102 707162 239546 707718
rect 240102 707162 275546 707718
rect 276102 707162 311546 707718
rect 312102 707162 347546 707718
rect 348102 707162 383546 707718
rect 384102 707162 419546 707718
rect 420102 707162 455546 707718
rect 456102 707162 491546 707718
rect 492102 707162 527546 707718
rect 528102 707162 563546 707718
rect 564102 707162 588222 707718
rect 588778 707162 588810 707718
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706202 -3894 706758
rect -3338 706202 5546 706758
rect 6102 706202 41546 706758
rect 42102 706202 77546 706758
rect 78102 706202 113546 706758
rect 114102 706202 149546 706758
rect 150102 706202 185546 706758
rect 186102 706202 221546 706758
rect 222102 706202 257546 706758
rect 258102 706202 293546 706758
rect 294102 706202 329546 706758
rect 330102 706202 365546 706758
rect 366102 706202 401546 706758
rect 402102 706202 437546 706758
rect 438102 706202 473546 706758
rect 474102 706202 509546 706758
rect 510102 706202 545546 706758
rect 546102 706202 581546 706758
rect 582102 706202 587262 706758
rect 587818 706202 587850 706758
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705242 -2934 705798
rect -2378 705242 19826 705798
rect 20382 705242 55826 705798
rect 56382 705242 91826 705798
rect 92382 705242 127826 705798
rect 128382 705242 163826 705798
rect 164382 705242 199826 705798
rect 200382 705242 235826 705798
rect 236382 705242 271826 705798
rect 272382 705242 307826 705798
rect 308382 705242 343826 705798
rect 344382 705242 379826 705798
rect 380382 705242 415826 705798
rect 416382 705242 451826 705798
rect 452382 705242 487826 705798
rect 488382 705242 523826 705798
rect 524382 705242 559826 705798
rect 560382 705242 586302 705798
rect 586858 705242 586890 705798
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704282 -1974 704838
rect -1418 704282 1826 704838
rect 2382 704282 37826 704838
rect 38382 704282 73826 704838
rect 74382 704282 109826 704838
rect 110382 704282 145826 704838
rect 146382 704282 181826 704838
rect 182382 704282 217826 704838
rect 218382 704282 253826 704838
rect 254382 704282 289826 704838
rect 290382 704282 325826 704838
rect 326382 704282 361826 704838
rect 362382 704282 397826 704838
rect 398382 704282 433826 704838
rect 434382 704282 469826 704838
rect 470382 704282 505826 704838
rect 506382 704282 541826 704838
rect 542382 704282 577826 704838
rect 578382 704282 585342 704838
rect 585898 704282 585930 704838
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698058 -7734 698614
rect -7178 698058 12986 698614
rect 13542 698058 48986 698614
rect 49542 698058 84986 698614
rect 85542 698058 120986 698614
rect 121542 698058 156986 698614
rect 157542 698058 192986 698614
rect 193542 698058 228986 698614
rect 229542 698058 264986 698614
rect 265542 698058 300986 698614
rect 301542 698058 336986 698614
rect 337542 698058 372986 698614
rect 373542 698058 408986 698614
rect 409542 698058 444986 698614
rect 445542 698058 480986 698614
rect 481542 698058 516986 698614
rect 517542 698058 552986 698614
rect 553542 698058 591102 698614
rect 591658 698058 592650 698614
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694338 -5814 694894
rect -5258 694338 9266 694894
rect 9822 694338 45266 694894
rect 45822 694338 81266 694894
rect 81822 694338 117266 694894
rect 117822 694338 153266 694894
rect 153822 694338 189266 694894
rect 189822 694338 225266 694894
rect 225822 694338 261266 694894
rect 261822 694338 297266 694894
rect 297822 694338 333266 694894
rect 333822 694338 369266 694894
rect 369822 694338 405266 694894
rect 405822 694338 441266 694894
rect 441822 694338 477266 694894
rect 477822 694338 513266 694894
rect 513822 694338 549266 694894
rect 549822 694338 589182 694894
rect 589738 694338 590730 694894
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690618 -3894 691174
rect -3338 690618 5546 691174
rect 6102 690618 41546 691174
rect 42102 690618 77546 691174
rect 78102 690618 113546 691174
rect 114102 690618 149546 691174
rect 150102 690618 185546 691174
rect 186102 690618 221546 691174
rect 222102 690618 257546 691174
rect 258102 690618 293546 691174
rect 294102 690618 329546 691174
rect 330102 690618 365546 691174
rect 366102 690618 401546 691174
rect 402102 690618 437546 691174
rect 438102 690618 473546 691174
rect 474102 690618 509546 691174
rect 510102 690618 545546 691174
rect 546102 690618 581546 691174
rect 582102 690618 587262 691174
rect 587818 690618 588810 691174
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 686898 -1974 687454
rect -1418 686898 1826 687454
rect 2382 686898 37826 687454
rect 38382 686898 73826 687454
rect 74382 686898 109826 687454
rect 110382 686898 145826 687454
rect 146382 686898 181826 687454
rect 182382 686898 217826 687454
rect 218382 686898 253826 687454
rect 254382 686898 289826 687454
rect 290382 686898 325826 687454
rect 326382 686898 361826 687454
rect 362382 686898 397826 687454
rect 398382 686898 433826 687454
rect 434382 686898 469826 687454
rect 470382 686898 505826 687454
rect 506382 686898 541826 687454
rect 542382 686898 577826 687454
rect 578382 686898 585342 687454
rect 585898 686898 586890 687454
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680058 -8694 680614
rect -8138 680058 30986 680614
rect 31542 680058 66986 680614
rect 67542 680058 102986 680614
rect 103542 680058 138986 680614
rect 139542 680058 174986 680614
rect 175542 680058 210986 680614
rect 211542 680058 246986 680614
rect 247542 680058 282986 680614
rect 283542 680058 318986 680614
rect 319542 680058 354986 680614
rect 355542 680058 390986 680614
rect 391542 680058 426986 680614
rect 427542 680058 462986 680614
rect 463542 680058 498986 680614
rect 499542 680058 534986 680614
rect 535542 680058 570986 680614
rect 571542 680058 592062 680614
rect 592618 680058 592650 680614
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676338 -6774 676894
rect -6218 676338 27266 676894
rect 27822 676338 63266 676894
rect 63822 676338 99266 676894
rect 99822 676338 135266 676894
rect 135822 676338 171266 676894
rect 171822 676338 207266 676894
rect 207822 676338 243266 676894
rect 243822 676338 279266 676894
rect 279822 676338 315266 676894
rect 315822 676338 351266 676894
rect 351822 676338 387266 676894
rect 387822 676338 423266 676894
rect 423822 676338 459266 676894
rect 459822 676338 495266 676894
rect 495822 676338 531266 676894
rect 531822 676338 567266 676894
rect 567822 676338 590142 676894
rect 590698 676338 590730 676894
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672618 -4854 673174
rect -4298 672618 23546 673174
rect 24102 672618 59546 673174
rect 60102 672618 95546 673174
rect 96102 672618 131546 673174
rect 132102 672618 167546 673174
rect 168102 672618 203546 673174
rect 204102 672618 239546 673174
rect 240102 672618 275546 673174
rect 276102 672618 311546 673174
rect 312102 672618 347546 673174
rect 348102 672618 383546 673174
rect 384102 672618 419546 673174
rect 420102 672618 455546 673174
rect 456102 672618 491546 673174
rect 492102 672618 527546 673174
rect 528102 672618 563546 673174
rect 564102 672618 588222 673174
rect 588778 672618 588810 673174
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 668898 -2934 669454
rect -2378 668898 19826 669454
rect 20382 668898 55826 669454
rect 56382 668898 91826 669454
rect 92382 668898 127826 669454
rect 128382 668898 163826 669454
rect 164382 668898 199826 669454
rect 200382 668898 235826 669454
rect 236382 668898 271826 669454
rect 272382 668898 307826 669454
rect 308382 668898 343826 669454
rect 344382 668898 379826 669454
rect 380382 668898 415826 669454
rect 416382 668898 451826 669454
rect 452382 668898 487826 669454
rect 488382 668898 523826 669454
rect 524382 668898 559826 669454
rect 560382 668898 586302 669454
rect 586858 668898 586890 669454
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662058 -7734 662614
rect -7178 662058 12986 662614
rect 13542 662058 48986 662614
rect 49542 662058 84986 662614
rect 85542 662058 120986 662614
rect 121542 662058 156986 662614
rect 157542 662058 192986 662614
rect 193542 662058 228986 662614
rect 229542 662058 264986 662614
rect 265542 662058 300986 662614
rect 301542 662058 336986 662614
rect 337542 662058 372986 662614
rect 373542 662058 408986 662614
rect 409542 662058 444986 662614
rect 445542 662058 480986 662614
rect 481542 662058 516986 662614
rect 517542 662058 552986 662614
rect 553542 662058 591102 662614
rect 591658 662058 592650 662614
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658338 -5814 658894
rect -5258 658338 9266 658894
rect 9822 658338 45266 658894
rect 45822 658338 81266 658894
rect 81822 658338 117266 658894
rect 117822 658338 153266 658894
rect 153822 658338 189266 658894
rect 189822 658338 225266 658894
rect 225822 658338 261266 658894
rect 261822 658338 297266 658894
rect 297822 658338 333266 658894
rect 333822 658338 369266 658894
rect 369822 658338 405266 658894
rect 405822 658338 441266 658894
rect 441822 658338 477266 658894
rect 477822 658338 513266 658894
rect 513822 658338 549266 658894
rect 549822 658338 589182 658894
rect 589738 658338 590730 658894
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654618 -3894 655174
rect -3338 654618 5546 655174
rect 6102 654618 41546 655174
rect 42102 654618 77546 655174
rect 78102 654618 113546 655174
rect 114102 654618 149546 655174
rect 150102 654618 185546 655174
rect 186102 654618 221546 655174
rect 222102 654618 257546 655174
rect 258102 654618 293546 655174
rect 294102 654618 329546 655174
rect 330102 654618 365546 655174
rect 366102 654618 401546 655174
rect 402102 654618 437546 655174
rect 438102 654618 473546 655174
rect 474102 654618 509546 655174
rect 510102 654618 545546 655174
rect 546102 654618 581546 655174
rect 582102 654618 587262 655174
rect 587818 654618 588810 655174
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 650898 -1974 651454
rect -1418 650898 1826 651454
rect 2382 650898 37826 651454
rect 38382 650898 73826 651454
rect 74382 650898 109826 651454
rect 110382 650898 145826 651454
rect 146382 650898 181826 651454
rect 182382 650898 217826 651454
rect 218382 650898 253826 651454
rect 254382 650898 289826 651454
rect 290382 650898 325826 651454
rect 326382 650898 361826 651454
rect 362382 650898 397826 651454
rect 398382 650898 433826 651454
rect 434382 650898 469826 651454
rect 470382 650898 505826 651454
rect 506382 650898 541826 651454
rect 542382 650898 577826 651454
rect 578382 650898 585342 651454
rect 585898 650898 586890 651454
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644058 -8694 644614
rect -8138 644058 30986 644614
rect 31542 644058 66986 644614
rect 67542 644058 102986 644614
rect 103542 644058 138986 644614
rect 139542 644058 174986 644614
rect 175542 644058 210986 644614
rect 211542 644058 246986 644614
rect 247542 644058 282986 644614
rect 283542 644058 318986 644614
rect 319542 644058 354986 644614
rect 355542 644058 390986 644614
rect 391542 644058 426986 644614
rect 427542 644058 462986 644614
rect 463542 644058 498986 644614
rect 499542 644058 534986 644614
rect 535542 644058 570986 644614
rect 571542 644058 592062 644614
rect 592618 644058 592650 644614
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640338 -6774 640894
rect -6218 640338 27266 640894
rect 27822 640338 63266 640894
rect 63822 640338 99266 640894
rect 99822 640338 135266 640894
rect 135822 640338 171266 640894
rect 171822 640338 207266 640894
rect 207822 640338 243266 640894
rect 243822 640338 279266 640894
rect 279822 640338 315266 640894
rect 315822 640338 351266 640894
rect 351822 640338 387266 640894
rect 387822 640338 423266 640894
rect 423822 640338 459266 640894
rect 459822 640338 495266 640894
rect 495822 640338 531266 640894
rect 531822 640338 567266 640894
rect 567822 640338 590142 640894
rect 590698 640338 590730 640894
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636618 -4854 637174
rect -4298 636618 23546 637174
rect 24102 636618 59546 637174
rect 60102 636618 95546 637174
rect 96102 636618 131546 637174
rect 132102 636618 167546 637174
rect 168102 636618 203546 637174
rect 204102 636618 239546 637174
rect 240102 636618 275546 637174
rect 276102 636618 311546 637174
rect 312102 636618 347546 637174
rect 348102 636618 383546 637174
rect 384102 636618 419546 637174
rect 420102 636618 455546 637174
rect 456102 636618 491546 637174
rect 492102 636618 527546 637174
rect 528102 636618 563546 637174
rect 564102 636618 588222 637174
rect 588778 636618 588810 637174
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 632898 -2934 633454
rect -2378 632898 19826 633454
rect 20382 632898 55826 633454
rect 56382 632898 91826 633454
rect 92382 632898 127826 633454
rect 128382 632898 163826 633454
rect 164382 632898 199826 633454
rect 200382 632898 235826 633454
rect 236382 632898 271826 633454
rect 272382 632898 307826 633454
rect 308382 632898 343826 633454
rect 344382 632898 379826 633454
rect 380382 632898 415826 633454
rect 416382 632898 451826 633454
rect 452382 632898 487826 633454
rect 488382 632898 523826 633454
rect 524382 632898 559826 633454
rect 560382 632898 586302 633454
rect 586858 632898 586890 633454
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626058 -7734 626614
rect -7178 626058 12986 626614
rect 13542 626058 48986 626614
rect 49542 626058 84986 626614
rect 85542 626058 120986 626614
rect 121542 626058 156986 626614
rect 157542 626058 192986 626614
rect 193542 626058 228986 626614
rect 229542 626058 264986 626614
rect 265542 626058 300986 626614
rect 301542 626058 336986 626614
rect 337542 626058 372986 626614
rect 373542 626058 408986 626614
rect 409542 626058 444986 626614
rect 445542 626058 480986 626614
rect 481542 626058 516986 626614
rect 517542 626058 552986 626614
rect 553542 626058 591102 626614
rect 591658 626058 592650 626614
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622338 -5814 622894
rect -5258 622338 9266 622894
rect 9822 622338 45266 622894
rect 45822 622338 81266 622894
rect 81822 622338 117266 622894
rect 117822 622338 153266 622894
rect 153822 622338 189266 622894
rect 189822 622338 225266 622894
rect 225822 622338 261266 622894
rect 261822 622338 297266 622894
rect 297822 622338 333266 622894
rect 333822 622338 369266 622894
rect 369822 622338 405266 622894
rect 405822 622338 441266 622894
rect 441822 622338 477266 622894
rect 477822 622338 513266 622894
rect 513822 622338 549266 622894
rect 549822 622338 589182 622894
rect 589738 622338 590730 622894
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618618 -3894 619174
rect -3338 618618 5546 619174
rect 6102 618618 41546 619174
rect 42102 618618 77546 619174
rect 78102 618618 113546 619174
rect 114102 618618 149546 619174
rect 150102 618618 185546 619174
rect 186102 618618 221546 619174
rect 222102 618618 257546 619174
rect 258102 618618 293546 619174
rect 294102 618618 329546 619174
rect 330102 618618 365546 619174
rect 366102 618618 401546 619174
rect 402102 618618 437546 619174
rect 438102 618618 473546 619174
rect 474102 618618 509546 619174
rect 510102 618618 545546 619174
rect 546102 618618 581546 619174
rect 582102 618618 587262 619174
rect 587818 618618 588810 619174
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 614898 -1974 615454
rect -1418 614898 1826 615454
rect 2382 614898 37826 615454
rect 38382 614898 73826 615454
rect 74382 614898 109826 615454
rect 110382 614898 145826 615454
rect 146382 614898 181826 615454
rect 182382 614898 217826 615454
rect 218382 614898 253826 615454
rect 254382 614898 289826 615454
rect 290382 614898 325826 615454
rect 326382 614898 361826 615454
rect 362382 614898 397826 615454
rect 398382 614898 433826 615454
rect 434382 614898 469826 615454
rect 470382 614898 505826 615454
rect 506382 614898 541826 615454
rect 542382 614898 577826 615454
rect 578382 614898 585342 615454
rect 585898 614898 586890 615454
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608058 -8694 608614
rect -8138 608058 30986 608614
rect 31542 608058 66986 608614
rect 67542 608058 102986 608614
rect 103542 608058 138986 608614
rect 139542 608058 174986 608614
rect 175542 608058 210986 608614
rect 211542 608058 246986 608614
rect 247542 608058 282986 608614
rect 283542 608058 318986 608614
rect 319542 608058 354986 608614
rect 355542 608058 390986 608614
rect 391542 608058 426986 608614
rect 427542 608058 462986 608614
rect 463542 608058 498986 608614
rect 499542 608058 534986 608614
rect 535542 608058 570986 608614
rect 571542 608058 592062 608614
rect 592618 608058 592650 608614
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604338 -6774 604894
rect -6218 604338 27266 604894
rect 27822 604338 63266 604894
rect 63822 604338 99266 604894
rect 99822 604338 135266 604894
rect 135822 604338 171266 604894
rect 171822 604338 207266 604894
rect 207822 604338 243266 604894
rect 243822 604338 279266 604894
rect 279822 604338 315266 604894
rect 315822 604338 351266 604894
rect 351822 604338 387266 604894
rect 387822 604338 423266 604894
rect 423822 604338 459266 604894
rect 459822 604338 495266 604894
rect 495822 604338 531266 604894
rect 531822 604338 567266 604894
rect 567822 604338 590142 604894
rect 590698 604338 590730 604894
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600618 -4854 601174
rect -4298 600618 23546 601174
rect 24102 600618 59546 601174
rect 60102 600618 95546 601174
rect 96102 600618 131546 601174
rect 132102 600618 167546 601174
rect 168102 600618 203546 601174
rect 204102 600618 239546 601174
rect 240102 600618 275546 601174
rect 276102 600618 311546 601174
rect 312102 600618 347546 601174
rect 348102 600618 383546 601174
rect 384102 600618 419546 601174
rect 420102 600618 455546 601174
rect 456102 600618 491546 601174
rect 492102 600618 527546 601174
rect 528102 600618 563546 601174
rect 564102 600618 588222 601174
rect 588778 600618 588810 601174
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 596898 -2934 597454
rect -2378 596898 19826 597454
rect 20382 596898 55826 597454
rect 56382 596898 91826 597454
rect 92382 596898 127826 597454
rect 128382 596898 163826 597454
rect 164382 596898 199826 597454
rect 200382 596898 235826 597454
rect 236382 596898 271826 597454
rect 272382 596898 307826 597454
rect 308382 596898 343826 597454
rect 344382 596898 379826 597454
rect 380382 596898 415826 597454
rect 416382 596898 451826 597454
rect 452382 596898 487826 597454
rect 488382 596898 523826 597454
rect 524382 596898 559826 597454
rect 560382 596898 586302 597454
rect 586858 596898 586890 597454
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590058 -7734 590614
rect -7178 590058 12986 590614
rect 13542 590058 48986 590614
rect 49542 590058 84986 590614
rect 85542 590058 120986 590614
rect 121542 590058 156986 590614
rect 157542 590058 192986 590614
rect 193542 590058 228986 590614
rect 229542 590058 264986 590614
rect 265542 590058 300986 590614
rect 301542 590058 336986 590614
rect 337542 590058 372986 590614
rect 373542 590058 408986 590614
rect 409542 590058 444986 590614
rect 445542 590058 480986 590614
rect 481542 590058 516986 590614
rect 517542 590058 552986 590614
rect 553542 590058 591102 590614
rect 591658 590058 592650 590614
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586338 -5814 586894
rect -5258 586338 9266 586894
rect 9822 586338 45266 586894
rect 45822 586338 81266 586894
rect 81822 586338 117266 586894
rect 117822 586338 153266 586894
rect 153822 586338 189266 586894
rect 189822 586338 225266 586894
rect 225822 586338 261266 586894
rect 261822 586338 297266 586894
rect 297822 586338 333266 586894
rect 333822 586338 369266 586894
rect 369822 586338 405266 586894
rect 405822 586338 441266 586894
rect 441822 586338 477266 586894
rect 477822 586338 513266 586894
rect 513822 586338 549266 586894
rect 549822 586338 589182 586894
rect 589738 586338 590730 586894
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582618 -3894 583174
rect -3338 582618 5546 583174
rect 6102 582618 41546 583174
rect 42102 582618 77546 583174
rect 78102 582618 113546 583174
rect 114102 582618 149546 583174
rect 150102 582618 185546 583174
rect 186102 582618 221546 583174
rect 222102 582618 257546 583174
rect 258102 582618 293546 583174
rect 294102 582618 329546 583174
rect 330102 582618 365546 583174
rect 366102 582618 401546 583174
rect 402102 582618 437546 583174
rect 438102 582618 473546 583174
rect 474102 582618 509546 583174
rect 510102 582618 545546 583174
rect 546102 582618 581546 583174
rect 582102 582618 587262 583174
rect 587818 582618 588810 583174
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 578898 -1974 579454
rect -1418 578898 1826 579454
rect 2382 578898 37826 579454
rect 38382 578898 73826 579454
rect 74382 578898 109826 579454
rect 110382 578898 145826 579454
rect 146382 578898 181826 579454
rect 182382 578898 217826 579454
rect 218382 578898 253826 579454
rect 254382 578898 289826 579454
rect 290382 578898 325826 579454
rect 326382 578898 361826 579454
rect 362382 578898 397826 579454
rect 398382 578898 433826 579454
rect 434382 578898 469826 579454
rect 470382 578898 505826 579454
rect 506382 578898 541826 579454
rect 542382 578898 577826 579454
rect 578382 578898 585342 579454
rect 585898 578898 586890 579454
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572058 -8694 572614
rect -8138 572058 30986 572614
rect 31542 572058 66986 572614
rect 67542 572058 102986 572614
rect 103542 572058 138986 572614
rect 139542 572058 174986 572614
rect 175542 572058 210986 572614
rect 211542 572058 246986 572614
rect 247542 572058 282986 572614
rect 283542 572058 318986 572614
rect 319542 572058 354986 572614
rect 355542 572058 390986 572614
rect 391542 572058 426986 572614
rect 427542 572058 462986 572614
rect 463542 572058 498986 572614
rect 499542 572058 534986 572614
rect 535542 572058 570986 572614
rect 571542 572058 592062 572614
rect 592618 572058 592650 572614
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568338 -6774 568894
rect -6218 568338 27266 568894
rect 27822 568338 63266 568894
rect 63822 568338 99266 568894
rect 99822 568338 135266 568894
rect 135822 568338 171266 568894
rect 171822 568338 207266 568894
rect 207822 568338 243266 568894
rect 243822 568338 279266 568894
rect 279822 568338 315266 568894
rect 315822 568338 351266 568894
rect 351822 568338 387266 568894
rect 387822 568338 423266 568894
rect 423822 568338 459266 568894
rect 459822 568338 495266 568894
rect 495822 568338 531266 568894
rect 531822 568338 567266 568894
rect 567822 568338 590142 568894
rect 590698 568338 590730 568894
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564618 -4854 565174
rect -4298 564618 23546 565174
rect 24102 564618 59546 565174
rect 60102 564618 95546 565174
rect 96102 564618 131546 565174
rect 132102 564618 167546 565174
rect 168102 564618 203546 565174
rect 204102 564618 239546 565174
rect 240102 564618 275546 565174
rect 276102 564618 311546 565174
rect 312102 564618 347546 565174
rect 348102 564618 383546 565174
rect 384102 564618 419546 565174
rect 420102 564618 455546 565174
rect 456102 564618 491546 565174
rect 492102 564618 527546 565174
rect 528102 564618 563546 565174
rect 564102 564618 588222 565174
rect 588778 564618 588810 565174
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 560898 -2934 561454
rect -2378 560898 19826 561454
rect 20382 560898 55826 561454
rect 56382 560898 91826 561454
rect 92382 560898 127826 561454
rect 128382 560898 163826 561454
rect 164382 560898 199826 561454
rect 200382 560898 235826 561454
rect 236382 560898 271826 561454
rect 272382 560898 307826 561454
rect 308382 560898 343826 561454
rect 344382 560898 379826 561454
rect 380382 560898 415826 561454
rect 416382 560898 451826 561454
rect 452382 560898 487826 561454
rect 488382 560898 523826 561454
rect 524382 560898 559826 561454
rect 560382 560898 586302 561454
rect 586858 560898 586890 561454
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554058 -7734 554614
rect -7178 554058 12986 554614
rect 13542 554058 48986 554614
rect 49542 554058 84986 554614
rect 85542 554058 120986 554614
rect 121542 554058 156986 554614
rect 157542 554058 192986 554614
rect 193542 554058 228986 554614
rect 229542 554058 264986 554614
rect 265542 554058 300986 554614
rect 301542 554058 336986 554614
rect 337542 554058 372986 554614
rect 373542 554058 408986 554614
rect 409542 554058 444986 554614
rect 445542 554058 480986 554614
rect 481542 554058 516986 554614
rect 517542 554058 552986 554614
rect 553542 554058 591102 554614
rect 591658 554058 592650 554614
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550338 -5814 550894
rect -5258 550338 9266 550894
rect 9822 550338 45266 550894
rect 45822 550338 81266 550894
rect 81822 550338 117266 550894
rect 117822 550338 153266 550894
rect 153822 550338 189266 550894
rect 189822 550338 225266 550894
rect 225822 550338 261266 550894
rect 261822 550338 297266 550894
rect 297822 550338 333266 550894
rect 333822 550338 369266 550894
rect 369822 550338 405266 550894
rect 405822 550338 441266 550894
rect 441822 550338 477266 550894
rect 477822 550338 513266 550894
rect 513822 550338 549266 550894
rect 549822 550338 589182 550894
rect 589738 550338 590730 550894
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546618 -3894 547174
rect -3338 546618 5546 547174
rect 6102 546618 41546 547174
rect 42102 546618 77546 547174
rect 78102 546618 113546 547174
rect 114102 546618 149546 547174
rect 150102 546618 185546 547174
rect 186102 546618 221546 547174
rect 222102 546618 257546 547174
rect 258102 546618 293546 547174
rect 294102 546618 329546 547174
rect 330102 546618 365546 547174
rect 366102 546618 401546 547174
rect 402102 546618 437546 547174
rect 438102 546618 473546 547174
rect 474102 546618 509546 547174
rect 510102 546618 545546 547174
rect 546102 546618 581546 547174
rect 582102 546618 587262 547174
rect 587818 546618 588810 547174
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 542898 -1974 543454
rect -1418 542898 1826 543454
rect 2382 542898 37826 543454
rect 38382 542898 73826 543454
rect 74382 542898 109826 543454
rect 110382 542898 145826 543454
rect 146382 542898 181826 543454
rect 182382 542898 217826 543454
rect 218382 542898 253826 543454
rect 254382 542898 289826 543454
rect 290382 542898 325826 543454
rect 326382 542898 361826 543454
rect 362382 542898 397826 543454
rect 398382 542898 433826 543454
rect 434382 542898 469826 543454
rect 470382 542898 505826 543454
rect 506382 542898 541826 543454
rect 542382 542898 577826 543454
rect 578382 542898 585342 543454
rect 585898 542898 586890 543454
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536058 -8694 536614
rect -8138 536058 30986 536614
rect 31542 536058 66986 536614
rect 67542 536058 102986 536614
rect 103542 536058 138986 536614
rect 139542 536058 174986 536614
rect 175542 536058 210986 536614
rect 211542 536058 246986 536614
rect 247542 536058 282986 536614
rect 283542 536058 318986 536614
rect 319542 536058 354986 536614
rect 355542 536058 390986 536614
rect 391542 536058 426986 536614
rect 427542 536058 462986 536614
rect 463542 536058 498986 536614
rect 499542 536058 534986 536614
rect 535542 536058 570986 536614
rect 571542 536058 592062 536614
rect 592618 536058 592650 536614
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532338 -6774 532894
rect -6218 532338 27266 532894
rect 27822 532338 63266 532894
rect 63822 532338 99266 532894
rect 99822 532338 135266 532894
rect 135822 532338 171266 532894
rect 171822 532338 207266 532894
rect 207822 532338 243266 532894
rect 243822 532338 279266 532894
rect 279822 532338 315266 532894
rect 315822 532338 351266 532894
rect 351822 532338 387266 532894
rect 387822 532338 423266 532894
rect 423822 532338 459266 532894
rect 459822 532338 495266 532894
rect 495822 532338 531266 532894
rect 531822 532338 567266 532894
rect 567822 532338 590142 532894
rect 590698 532338 590730 532894
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528618 -4854 529174
rect -4298 528618 23546 529174
rect 24102 528618 59546 529174
rect 60102 528618 95546 529174
rect 96102 528618 131546 529174
rect 132102 528618 167546 529174
rect 168102 528618 203546 529174
rect 204102 528618 239546 529174
rect 240102 528618 275546 529174
rect 276102 528618 311546 529174
rect 312102 528618 347546 529174
rect 348102 528618 383546 529174
rect 384102 528618 419546 529174
rect 420102 528618 455546 529174
rect 456102 528618 491546 529174
rect 492102 528618 527546 529174
rect 528102 528618 563546 529174
rect 564102 528618 588222 529174
rect 588778 528618 588810 529174
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 524898 -2934 525454
rect -2378 524898 19826 525454
rect 20382 524898 55826 525454
rect 56382 524898 91826 525454
rect 92382 524898 127826 525454
rect 128382 524898 163826 525454
rect 164382 524898 199826 525454
rect 200382 524898 235826 525454
rect 236382 524898 271826 525454
rect 272382 524898 307826 525454
rect 308382 524898 343826 525454
rect 344382 524898 379826 525454
rect 380382 524898 415826 525454
rect 416382 524898 451826 525454
rect 452382 524898 487826 525454
rect 488382 524898 523826 525454
rect 524382 524898 559826 525454
rect 560382 524898 586302 525454
rect 586858 524898 586890 525454
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518058 -7734 518614
rect -7178 518058 12986 518614
rect 13542 518058 48986 518614
rect 49542 518058 84986 518614
rect 85542 518058 120986 518614
rect 121542 518058 156986 518614
rect 157542 518058 192986 518614
rect 193542 518058 228986 518614
rect 229542 518058 264986 518614
rect 265542 518058 300986 518614
rect 301542 518058 336986 518614
rect 337542 518058 372986 518614
rect 373542 518058 408986 518614
rect 409542 518058 444986 518614
rect 445542 518058 480986 518614
rect 481542 518058 516986 518614
rect 517542 518058 552986 518614
rect 553542 518058 591102 518614
rect 591658 518058 592650 518614
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514338 -5814 514894
rect -5258 514338 9266 514894
rect 9822 514338 45266 514894
rect 45822 514338 81266 514894
rect 81822 514338 117266 514894
rect 117822 514338 153266 514894
rect 153822 514338 189266 514894
rect 189822 514338 225266 514894
rect 225822 514338 261266 514894
rect 261822 514338 297266 514894
rect 297822 514338 333266 514894
rect 333822 514338 369266 514894
rect 369822 514338 405266 514894
rect 405822 514338 441266 514894
rect 441822 514338 477266 514894
rect 477822 514338 513266 514894
rect 513822 514338 549266 514894
rect 549822 514338 589182 514894
rect 589738 514338 590730 514894
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510618 -3894 511174
rect -3338 510618 5546 511174
rect 6102 510618 41546 511174
rect 42102 510618 77546 511174
rect 78102 510618 113546 511174
rect 114102 510618 149546 511174
rect 150102 510618 185546 511174
rect 186102 510618 221546 511174
rect 222102 510618 257546 511174
rect 258102 510618 293546 511174
rect 294102 510618 329546 511174
rect 330102 510618 365546 511174
rect 366102 510618 401546 511174
rect 402102 510618 437546 511174
rect 438102 510618 473546 511174
rect 474102 510618 509546 511174
rect 510102 510618 545546 511174
rect 546102 510618 581546 511174
rect 582102 510618 587262 511174
rect 587818 510618 588810 511174
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 506898 -1974 507454
rect -1418 506898 1826 507454
rect 2382 506898 37826 507454
rect 38382 506898 73826 507454
rect 74382 506898 109826 507454
rect 110382 506898 145826 507454
rect 146382 506898 181826 507454
rect 182382 506898 217826 507454
rect 218382 506898 253826 507454
rect 254382 506898 289826 507454
rect 290382 506898 325826 507454
rect 326382 506898 361826 507454
rect 362382 506898 397826 507454
rect 398382 506898 433826 507454
rect 434382 506898 469826 507454
rect 470382 506898 505826 507454
rect 506382 506898 541826 507454
rect 542382 506898 577826 507454
rect 578382 506898 585342 507454
rect 585898 506898 586890 507454
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500058 -8694 500614
rect -8138 500058 30986 500614
rect 31542 500058 66986 500614
rect 67542 500058 102986 500614
rect 103542 500058 138986 500614
rect 139542 500058 174986 500614
rect 175542 500058 210986 500614
rect 211542 500058 246986 500614
rect 247542 500058 282986 500614
rect 283542 500058 318986 500614
rect 319542 500058 354986 500614
rect 355542 500058 390986 500614
rect 391542 500058 426986 500614
rect 427542 500058 462986 500614
rect 463542 500058 498986 500614
rect 499542 500058 534986 500614
rect 535542 500058 570986 500614
rect 571542 500058 592062 500614
rect 592618 500058 592650 500614
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496338 -6774 496894
rect -6218 496338 27266 496894
rect 27822 496338 63266 496894
rect 63822 496338 99266 496894
rect 99822 496338 135266 496894
rect 135822 496338 171266 496894
rect 171822 496338 207266 496894
rect 207822 496338 243266 496894
rect 243822 496338 279266 496894
rect 279822 496338 315266 496894
rect 315822 496338 351266 496894
rect 351822 496338 387266 496894
rect 387822 496338 423266 496894
rect 423822 496338 459266 496894
rect 459822 496338 495266 496894
rect 495822 496338 531266 496894
rect 531822 496338 567266 496894
rect 567822 496338 590142 496894
rect 590698 496338 590730 496894
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492618 -4854 493174
rect -4298 492618 23546 493174
rect 24102 492618 59546 493174
rect 60102 492618 95546 493174
rect 96102 492618 131546 493174
rect 132102 492618 167546 493174
rect 168102 492618 203546 493174
rect 204102 492618 239546 493174
rect 240102 492618 275546 493174
rect 276102 492618 311546 493174
rect 312102 492618 347546 493174
rect 348102 492618 383546 493174
rect 384102 492618 419546 493174
rect 420102 492618 455546 493174
rect 456102 492618 491546 493174
rect 492102 492618 527546 493174
rect 528102 492618 563546 493174
rect 564102 492618 588222 493174
rect 588778 492618 588810 493174
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 488898 -2934 489454
rect -2378 488898 19826 489454
rect 20382 488898 55826 489454
rect 56382 488898 91826 489454
rect 92382 488898 127826 489454
rect 128382 488898 163826 489454
rect 164382 488898 199826 489454
rect 200382 488898 235826 489454
rect 236382 488898 271826 489454
rect 272382 488898 307826 489454
rect 308382 488898 343826 489454
rect 344382 488898 379826 489454
rect 380382 488898 415826 489454
rect 416382 488898 451826 489454
rect 452382 488898 487826 489454
rect 488382 488898 523826 489454
rect 524382 488898 559826 489454
rect 560382 488898 586302 489454
rect 586858 488898 586890 489454
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482058 -7734 482614
rect -7178 482058 12986 482614
rect 13542 482058 48986 482614
rect 49542 482058 84986 482614
rect 85542 482058 120986 482614
rect 121542 482058 156986 482614
rect 157542 482058 192986 482614
rect 193542 482058 228986 482614
rect 229542 482058 264986 482614
rect 265542 482058 300986 482614
rect 301542 482058 336986 482614
rect 337542 482058 372986 482614
rect 373542 482058 408986 482614
rect 409542 482058 444986 482614
rect 445542 482058 480986 482614
rect 481542 482058 516986 482614
rect 517542 482058 552986 482614
rect 553542 482058 591102 482614
rect 591658 482058 592650 482614
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478338 -5814 478894
rect -5258 478338 9266 478894
rect 9822 478338 45266 478894
rect 45822 478338 81266 478894
rect 81822 478338 117266 478894
rect 117822 478338 153266 478894
rect 153822 478338 189266 478894
rect 189822 478338 225266 478894
rect 225822 478338 261266 478894
rect 261822 478338 297266 478894
rect 297822 478338 333266 478894
rect 333822 478338 369266 478894
rect 369822 478338 405266 478894
rect 405822 478338 441266 478894
rect 441822 478338 477266 478894
rect 477822 478338 513266 478894
rect 513822 478338 549266 478894
rect 549822 478338 589182 478894
rect 589738 478338 590730 478894
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474618 -3894 475174
rect -3338 474618 5546 475174
rect 6102 474618 41546 475174
rect 42102 474618 77546 475174
rect 78102 474618 113546 475174
rect 114102 474618 149546 475174
rect 150102 474618 185546 475174
rect 186102 474618 221546 475174
rect 222102 474618 257546 475174
rect 258102 474618 293546 475174
rect 294102 474618 329546 475174
rect 330102 474618 365546 475174
rect 366102 474618 401546 475174
rect 402102 474618 437546 475174
rect 438102 474618 473546 475174
rect 474102 474618 509546 475174
rect 510102 474618 545546 475174
rect 546102 474618 581546 475174
rect 582102 474618 587262 475174
rect 587818 474618 588810 475174
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 470898 -1974 471454
rect -1418 470898 1826 471454
rect 2382 470898 37826 471454
rect 38382 470898 73826 471454
rect 74382 470898 109826 471454
rect 110382 470898 145826 471454
rect 146382 470898 181826 471454
rect 182382 470898 217826 471454
rect 218382 470898 253826 471454
rect 254382 470898 289826 471454
rect 290382 470898 325826 471454
rect 326382 470898 361826 471454
rect 362382 470898 397826 471454
rect 398382 470898 433826 471454
rect 434382 470898 469826 471454
rect 470382 470898 505826 471454
rect 506382 470898 541826 471454
rect 542382 470898 577826 471454
rect 578382 470898 585342 471454
rect 585898 470898 586890 471454
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464058 -8694 464614
rect -8138 464058 30986 464614
rect 31542 464058 66986 464614
rect 67542 464058 102986 464614
rect 103542 464058 138986 464614
rect 139542 464058 174986 464614
rect 175542 464058 210986 464614
rect 211542 464058 246986 464614
rect 247542 464058 282986 464614
rect 283542 464058 318986 464614
rect 319542 464058 354986 464614
rect 355542 464058 390986 464614
rect 391542 464058 426986 464614
rect 427542 464058 462986 464614
rect 463542 464058 498986 464614
rect 499542 464058 534986 464614
rect 535542 464058 570986 464614
rect 571542 464058 592062 464614
rect 592618 464058 592650 464614
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460338 -6774 460894
rect -6218 460338 27266 460894
rect 27822 460338 63266 460894
rect 63822 460338 99266 460894
rect 99822 460338 135266 460894
rect 135822 460338 171266 460894
rect 171822 460338 207266 460894
rect 207822 460338 243266 460894
rect 243822 460338 279266 460894
rect 279822 460338 315266 460894
rect 315822 460338 351266 460894
rect 351822 460338 387266 460894
rect 387822 460338 423266 460894
rect 423822 460338 459266 460894
rect 459822 460338 495266 460894
rect 495822 460338 531266 460894
rect 531822 460338 567266 460894
rect 567822 460338 590142 460894
rect 590698 460338 590730 460894
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456618 -4854 457174
rect -4298 456618 23546 457174
rect 24102 456618 59546 457174
rect 60102 456618 95546 457174
rect 96102 456618 131546 457174
rect 132102 456618 167546 457174
rect 168102 456618 203546 457174
rect 204102 456618 419546 457174
rect 420102 456618 455546 457174
rect 456102 456618 491546 457174
rect 492102 456618 527546 457174
rect 528102 456618 563546 457174
rect 564102 456618 588222 457174
rect 588778 456618 588810 457174
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 452898 -2934 453454
rect -2378 452898 19826 453454
rect 20382 452898 55826 453454
rect 56382 452898 91826 453454
rect 92382 452898 127826 453454
rect 128382 452898 163826 453454
rect 164382 452898 199826 453454
rect 200382 453218 254610 453454
rect 254846 453218 285330 453454
rect 285566 453218 316050 453454
rect 316286 453218 346770 453454
rect 347006 453218 377490 453454
rect 377726 453218 408210 453454
rect 408446 453218 415826 453454
rect 200382 453134 415826 453218
rect 200382 452898 254610 453134
rect 254846 452898 285330 453134
rect 285566 452898 316050 453134
rect 316286 452898 346770 453134
rect 347006 452898 377490 453134
rect 377726 452898 408210 453134
rect 408446 452898 415826 453134
rect 416382 452898 451826 453454
rect 452382 452898 487826 453454
rect 488382 452898 523826 453454
rect 524382 452898 559826 453454
rect 560382 452898 586302 453454
rect 586858 452898 586890 453454
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446058 -7734 446614
rect -7178 446058 12986 446614
rect 13542 446058 48986 446614
rect 49542 446058 84986 446614
rect 85542 446058 120986 446614
rect 121542 446058 156986 446614
rect 157542 446058 192986 446614
rect 193542 446058 228986 446614
rect 229542 446058 444986 446614
rect 445542 446058 480986 446614
rect 481542 446058 516986 446614
rect 517542 446058 552986 446614
rect 553542 446058 591102 446614
rect 591658 446058 592650 446614
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442338 -5814 442894
rect -5258 442338 9266 442894
rect 9822 442338 45266 442894
rect 45822 442338 81266 442894
rect 81822 442338 117266 442894
rect 117822 442338 153266 442894
rect 153822 442338 189266 442894
rect 189822 442338 225266 442894
rect 225822 442338 441266 442894
rect 441822 442338 477266 442894
rect 477822 442338 513266 442894
rect 513822 442338 549266 442894
rect 549822 442338 589182 442894
rect 589738 442338 590730 442894
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438618 -3894 439174
rect -3338 438618 5546 439174
rect 6102 438618 41546 439174
rect 42102 438618 77546 439174
rect 78102 438618 113546 439174
rect 114102 438618 149546 439174
rect 150102 438618 185546 439174
rect 186102 438618 221546 439174
rect 222102 438618 437546 439174
rect 438102 438618 473546 439174
rect 474102 438618 509546 439174
rect 510102 438618 545546 439174
rect 546102 438618 581546 439174
rect 582102 438618 587262 439174
rect 587818 438618 588810 439174
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 434898 -1974 435454
rect -1418 434898 1826 435454
rect 2382 434898 37826 435454
rect 38382 434898 73826 435454
rect 74382 434898 109826 435454
rect 110382 434898 145826 435454
rect 146382 434898 181826 435454
rect 182382 434898 217826 435454
rect 218382 435218 239250 435454
rect 239486 435218 269970 435454
rect 270206 435218 300690 435454
rect 300926 435218 331410 435454
rect 331646 435218 362130 435454
rect 362366 435218 392850 435454
rect 393086 435218 433826 435454
rect 218382 435134 433826 435218
rect 218382 434898 239250 435134
rect 239486 434898 269970 435134
rect 270206 434898 300690 435134
rect 300926 434898 331410 435134
rect 331646 434898 362130 435134
rect 362366 434898 392850 435134
rect 393086 434898 433826 435134
rect 434382 434898 469826 435454
rect 470382 434898 505826 435454
rect 506382 434898 541826 435454
rect 542382 434898 577826 435454
rect 578382 434898 585342 435454
rect 585898 434898 586890 435454
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428058 -8694 428614
rect -8138 428058 30986 428614
rect 31542 428058 66986 428614
rect 67542 428058 102986 428614
rect 103542 428058 138986 428614
rect 139542 428058 174986 428614
rect 175542 428058 210986 428614
rect 211542 428058 426986 428614
rect 427542 428058 462986 428614
rect 463542 428058 498986 428614
rect 499542 428058 534986 428614
rect 535542 428058 570986 428614
rect 571542 428058 592062 428614
rect 592618 428058 592650 428614
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424338 -6774 424894
rect -6218 424338 27266 424894
rect 27822 424338 63266 424894
rect 63822 424338 99266 424894
rect 99822 424338 135266 424894
rect 135822 424338 171266 424894
rect 171822 424338 207266 424894
rect 207822 424338 423266 424894
rect 423822 424338 459266 424894
rect 459822 424338 495266 424894
rect 495822 424338 531266 424894
rect 531822 424338 567266 424894
rect 567822 424338 590142 424894
rect 590698 424338 590730 424894
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420618 -4854 421174
rect -4298 420618 23546 421174
rect 24102 420618 59546 421174
rect 60102 420618 95546 421174
rect 96102 420618 131546 421174
rect 132102 420618 167546 421174
rect 168102 420618 203546 421174
rect 204102 420618 419546 421174
rect 420102 420618 455546 421174
rect 456102 420618 491546 421174
rect 492102 420618 527546 421174
rect 528102 420618 563546 421174
rect 564102 420618 588222 421174
rect 588778 420618 588810 421174
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 416898 -2934 417454
rect -2378 416898 19826 417454
rect 20382 416898 55826 417454
rect 56382 416898 91826 417454
rect 92382 416898 127826 417454
rect 128382 416898 163826 417454
rect 164382 416898 199826 417454
rect 200382 417218 254610 417454
rect 254846 417218 285330 417454
rect 285566 417218 316050 417454
rect 316286 417218 346770 417454
rect 347006 417218 377490 417454
rect 377726 417218 408210 417454
rect 408446 417218 415826 417454
rect 200382 417134 415826 417218
rect 200382 416898 254610 417134
rect 254846 416898 285330 417134
rect 285566 416898 316050 417134
rect 316286 416898 346770 417134
rect 347006 416898 377490 417134
rect 377726 416898 408210 417134
rect 408446 416898 415826 417134
rect 416382 416898 451826 417454
rect 452382 416898 487826 417454
rect 488382 416898 523826 417454
rect 524382 416898 559826 417454
rect 560382 416898 586302 417454
rect 586858 416898 586890 417454
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410058 -7734 410614
rect -7178 410058 12986 410614
rect 13542 410058 48986 410614
rect 49542 410058 84986 410614
rect 85542 410058 120986 410614
rect 121542 410058 156986 410614
rect 157542 410058 192986 410614
rect 193542 410058 228986 410614
rect 229542 410058 444986 410614
rect 445542 410058 480986 410614
rect 481542 410058 516986 410614
rect 517542 410058 552986 410614
rect 553542 410058 591102 410614
rect 591658 410058 592650 410614
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406338 -5814 406894
rect -5258 406338 9266 406894
rect 9822 406338 45266 406894
rect 45822 406338 81266 406894
rect 81822 406338 117266 406894
rect 117822 406338 153266 406894
rect 153822 406338 189266 406894
rect 189822 406338 225266 406894
rect 225822 406338 441266 406894
rect 441822 406338 477266 406894
rect 477822 406338 513266 406894
rect 513822 406338 549266 406894
rect 549822 406338 589182 406894
rect 589738 406338 590730 406894
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402618 -3894 403174
rect -3338 402618 5546 403174
rect 6102 402618 41546 403174
rect 42102 402618 77546 403174
rect 78102 402618 113546 403174
rect 114102 402618 149546 403174
rect 150102 402618 185546 403174
rect 186102 402618 221546 403174
rect 222102 402618 437546 403174
rect 438102 402618 473546 403174
rect 474102 402618 509546 403174
rect 510102 402618 545546 403174
rect 546102 402618 581546 403174
rect 582102 402618 587262 403174
rect 587818 402618 588810 403174
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 398898 -1974 399454
rect -1418 398898 1826 399454
rect 2382 398898 37826 399454
rect 38382 398898 73826 399454
rect 74382 398898 109826 399454
rect 110382 398898 145826 399454
rect 146382 398898 181826 399454
rect 182382 398898 217826 399454
rect 218382 399218 239250 399454
rect 239486 399218 269970 399454
rect 270206 399218 300690 399454
rect 300926 399218 331410 399454
rect 331646 399218 362130 399454
rect 362366 399218 392850 399454
rect 393086 399218 433826 399454
rect 218382 399134 433826 399218
rect 218382 398898 239250 399134
rect 239486 398898 269970 399134
rect 270206 398898 300690 399134
rect 300926 398898 331410 399134
rect 331646 398898 362130 399134
rect 362366 398898 392850 399134
rect 393086 398898 433826 399134
rect 434382 398898 469826 399454
rect 470382 398898 505826 399454
rect 506382 398898 541826 399454
rect 542382 398898 577826 399454
rect 578382 398898 585342 399454
rect 585898 398898 586890 399454
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392058 -8694 392614
rect -8138 392058 30986 392614
rect 31542 392058 66986 392614
rect 67542 392058 102986 392614
rect 103542 392058 138986 392614
rect 139542 392058 174986 392614
rect 175542 392058 210986 392614
rect 211542 392058 426986 392614
rect 427542 392058 462986 392614
rect 463542 392058 498986 392614
rect 499542 392058 534986 392614
rect 535542 392058 570986 392614
rect 571542 392058 592062 392614
rect 592618 392058 592650 392614
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388338 -6774 388894
rect -6218 388338 27266 388894
rect 27822 388338 63266 388894
rect 63822 388338 99266 388894
rect 99822 388338 135266 388894
rect 135822 388338 171266 388894
rect 171822 388338 207266 388894
rect 207822 388338 423266 388894
rect 423822 388338 459266 388894
rect 459822 388338 495266 388894
rect 495822 388338 531266 388894
rect 531822 388338 567266 388894
rect 567822 388338 590142 388894
rect 590698 388338 590730 388894
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384618 -4854 385174
rect -4298 384618 23546 385174
rect 24102 384618 59546 385174
rect 60102 384618 95546 385174
rect 96102 384618 131546 385174
rect 132102 384618 167546 385174
rect 168102 384618 203546 385174
rect 204102 384618 419546 385174
rect 420102 384618 455546 385174
rect 456102 384618 491546 385174
rect 492102 384618 527546 385174
rect 528102 384618 563546 385174
rect 564102 384618 588222 385174
rect 588778 384618 588810 385174
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 380898 -2934 381454
rect -2378 380898 19826 381454
rect 20382 380898 55826 381454
rect 56382 380898 91826 381454
rect 92382 380898 127826 381454
rect 128382 380898 163826 381454
rect 164382 380898 199826 381454
rect 200382 381218 254610 381454
rect 254846 381218 285330 381454
rect 285566 381218 316050 381454
rect 316286 381218 346770 381454
rect 347006 381218 377490 381454
rect 377726 381218 408210 381454
rect 408446 381218 415826 381454
rect 200382 381134 415826 381218
rect 200382 380898 254610 381134
rect 254846 380898 285330 381134
rect 285566 380898 316050 381134
rect 316286 380898 346770 381134
rect 347006 380898 377490 381134
rect 377726 380898 408210 381134
rect 408446 380898 415826 381134
rect 416382 380898 451826 381454
rect 452382 380898 487826 381454
rect 488382 380898 523826 381454
rect 524382 380898 559826 381454
rect 560382 380898 586302 381454
rect 586858 380898 586890 381454
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374058 -7734 374614
rect -7178 374058 12986 374614
rect 13542 374058 48986 374614
rect 49542 374058 84986 374614
rect 85542 374058 120986 374614
rect 121542 374058 156986 374614
rect 157542 374058 192986 374614
rect 193542 374058 228986 374614
rect 229542 374058 444986 374614
rect 445542 374058 480986 374614
rect 481542 374058 516986 374614
rect 517542 374058 552986 374614
rect 553542 374058 591102 374614
rect 591658 374058 592650 374614
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370338 -5814 370894
rect -5258 370338 9266 370894
rect 9822 370338 45266 370894
rect 45822 370338 81266 370894
rect 81822 370338 117266 370894
rect 117822 370338 153266 370894
rect 153822 370338 189266 370894
rect 189822 370338 225266 370894
rect 225822 370338 441266 370894
rect 441822 370338 477266 370894
rect 477822 370338 513266 370894
rect 513822 370338 549266 370894
rect 549822 370338 589182 370894
rect 589738 370338 590730 370894
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366618 -3894 367174
rect -3338 366618 5546 367174
rect 6102 366618 41546 367174
rect 42102 366618 77546 367174
rect 78102 366618 113546 367174
rect 114102 366618 149546 367174
rect 150102 366618 185546 367174
rect 186102 366618 221546 367174
rect 222102 366618 437546 367174
rect 438102 366618 473546 367174
rect 474102 366618 509546 367174
rect 510102 366618 545546 367174
rect 546102 366618 581546 367174
rect 582102 366618 587262 367174
rect 587818 366618 588810 367174
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 362898 -1974 363454
rect -1418 362898 1826 363454
rect 2382 362898 37826 363454
rect 38382 362898 73826 363454
rect 74382 362898 109826 363454
rect 110382 362898 145826 363454
rect 146382 362898 181826 363454
rect 182382 362898 217826 363454
rect 218382 363218 239250 363454
rect 239486 363218 269970 363454
rect 270206 363218 300690 363454
rect 300926 363218 331410 363454
rect 331646 363218 362130 363454
rect 362366 363218 392850 363454
rect 393086 363218 433826 363454
rect 218382 363134 433826 363218
rect 218382 362898 239250 363134
rect 239486 362898 269970 363134
rect 270206 362898 300690 363134
rect 300926 362898 331410 363134
rect 331646 362898 362130 363134
rect 362366 362898 392850 363134
rect 393086 362898 433826 363134
rect 434382 362898 469826 363454
rect 470382 362898 505826 363454
rect 506382 362898 541826 363454
rect 542382 362898 577826 363454
rect 578382 362898 585342 363454
rect 585898 362898 586890 363454
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356058 -8694 356614
rect -8138 356058 30986 356614
rect 31542 356058 66986 356614
rect 67542 356058 102986 356614
rect 103542 356058 138986 356614
rect 139542 356058 174986 356614
rect 175542 356058 210986 356614
rect 211542 356058 426986 356614
rect 427542 356058 462986 356614
rect 463542 356058 498986 356614
rect 499542 356058 534986 356614
rect 535542 356058 570986 356614
rect 571542 356058 592062 356614
rect 592618 356058 592650 356614
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352338 -6774 352894
rect -6218 352338 27266 352894
rect 27822 352338 63266 352894
rect 63822 352338 99266 352894
rect 99822 352338 135266 352894
rect 135822 352338 171266 352894
rect 171822 352338 207266 352894
rect 207822 352338 423266 352894
rect 423822 352338 459266 352894
rect 459822 352338 495266 352894
rect 495822 352338 531266 352894
rect 531822 352338 567266 352894
rect 567822 352338 590142 352894
rect 590698 352338 590730 352894
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348618 -4854 349174
rect -4298 348618 23546 349174
rect 24102 348618 59546 349174
rect 60102 348618 95546 349174
rect 96102 348618 131546 349174
rect 132102 348618 167546 349174
rect 168102 348618 203546 349174
rect 204102 348618 419546 349174
rect 420102 348618 455546 349174
rect 456102 348618 491546 349174
rect 492102 348618 527546 349174
rect 528102 348618 563546 349174
rect 564102 348618 588222 349174
rect 588778 348618 588810 349174
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 344898 -2934 345454
rect -2378 344898 19826 345454
rect 20382 344898 55826 345454
rect 56382 344898 91826 345454
rect 92382 344898 127826 345454
rect 128382 344898 163826 345454
rect 164382 344898 199826 345454
rect 200382 345218 254610 345454
rect 254846 345218 285330 345454
rect 285566 345218 316050 345454
rect 316286 345218 346770 345454
rect 347006 345218 377490 345454
rect 377726 345218 408210 345454
rect 408446 345218 415826 345454
rect 200382 345134 415826 345218
rect 200382 344898 254610 345134
rect 254846 344898 285330 345134
rect 285566 344898 316050 345134
rect 316286 344898 346770 345134
rect 347006 344898 377490 345134
rect 377726 344898 408210 345134
rect 408446 344898 415826 345134
rect 416382 344898 451826 345454
rect 452382 344898 487826 345454
rect 488382 344898 523826 345454
rect 524382 344898 559826 345454
rect 560382 344898 586302 345454
rect 586858 344898 586890 345454
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338058 -7734 338614
rect -7178 338058 12986 338614
rect 13542 338058 48986 338614
rect 49542 338058 84986 338614
rect 85542 338058 120986 338614
rect 121542 338058 156986 338614
rect 157542 338058 192986 338614
rect 193542 338058 228986 338614
rect 229542 338058 444986 338614
rect 445542 338058 480986 338614
rect 481542 338058 516986 338614
rect 517542 338058 552986 338614
rect 553542 338058 591102 338614
rect 591658 338058 592650 338614
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334338 -5814 334894
rect -5258 334338 9266 334894
rect 9822 334338 45266 334894
rect 45822 334338 81266 334894
rect 81822 334338 117266 334894
rect 117822 334338 153266 334894
rect 153822 334338 189266 334894
rect 189822 334338 225266 334894
rect 225822 334338 261266 334894
rect 261822 334338 297266 334894
rect 297822 334338 333266 334894
rect 333822 334338 369266 334894
rect 369822 334338 405266 334894
rect 405822 334338 441266 334894
rect 441822 334338 477266 334894
rect 477822 334338 513266 334894
rect 513822 334338 549266 334894
rect 549822 334338 589182 334894
rect 589738 334338 590730 334894
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330618 -3894 331174
rect -3338 330618 5546 331174
rect 6102 330618 41546 331174
rect 42102 330618 77546 331174
rect 78102 330618 113546 331174
rect 114102 330618 149546 331174
rect 150102 330618 185546 331174
rect 186102 330618 221546 331174
rect 222102 330618 257546 331174
rect 258102 330618 293546 331174
rect 294102 330618 329546 331174
rect 330102 330618 365546 331174
rect 366102 330618 401546 331174
rect 402102 330618 437546 331174
rect 438102 330618 473546 331174
rect 474102 330618 509546 331174
rect 510102 330618 545546 331174
rect 546102 330618 581546 331174
rect 582102 330618 587262 331174
rect 587818 330618 588810 331174
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 326898 -1974 327454
rect -1418 326898 1826 327454
rect 2382 326898 37826 327454
rect 38382 326898 73826 327454
rect 74382 326898 109826 327454
rect 110382 326898 145826 327454
rect 146382 326898 181826 327454
rect 182382 326898 217826 327454
rect 218382 326898 253826 327454
rect 254382 326898 289826 327454
rect 290382 326898 325826 327454
rect 326382 326898 361826 327454
rect 362382 326898 397826 327454
rect 398382 326898 433826 327454
rect 434382 326898 469826 327454
rect 470382 326898 505826 327454
rect 506382 326898 541826 327454
rect 542382 326898 577826 327454
rect 578382 326898 585342 327454
rect 585898 326898 586890 327454
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320058 -8694 320614
rect -8138 320058 30986 320614
rect 31542 320058 66986 320614
rect 67542 320058 102986 320614
rect 103542 320058 138986 320614
rect 139542 320058 174986 320614
rect 175542 320058 210986 320614
rect 211542 320058 246986 320614
rect 247542 320058 282986 320614
rect 283542 320058 318986 320614
rect 319542 320058 354986 320614
rect 355542 320058 390986 320614
rect 391542 320058 426986 320614
rect 427542 320058 462986 320614
rect 463542 320058 498986 320614
rect 499542 320058 534986 320614
rect 535542 320058 570986 320614
rect 571542 320058 592062 320614
rect 592618 320058 592650 320614
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316338 -6774 316894
rect -6218 316338 27266 316894
rect 27822 316338 63266 316894
rect 63822 316338 99266 316894
rect 99822 316338 135266 316894
rect 135822 316338 171266 316894
rect 171822 316338 207266 316894
rect 207822 316338 243266 316894
rect 243822 316338 279266 316894
rect 279822 316338 315266 316894
rect 315822 316338 351266 316894
rect 351822 316338 387266 316894
rect 387822 316338 423266 316894
rect 423822 316338 459266 316894
rect 459822 316338 495266 316894
rect 495822 316338 531266 316894
rect 531822 316338 567266 316894
rect 567822 316338 590142 316894
rect 590698 316338 590730 316894
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312618 -4854 313174
rect -4298 312618 23546 313174
rect 24102 312618 59546 313174
rect 60102 312618 95546 313174
rect 96102 312618 131546 313174
rect 132102 312618 167546 313174
rect 168102 312618 203546 313174
rect 204102 312618 239546 313174
rect 240102 312618 275546 313174
rect 276102 312618 311546 313174
rect 312102 312618 347546 313174
rect 348102 312618 383546 313174
rect 384102 312618 419546 313174
rect 420102 312618 455546 313174
rect 456102 312618 491546 313174
rect 492102 312618 527546 313174
rect 528102 312618 563546 313174
rect 564102 312618 588222 313174
rect 588778 312618 588810 313174
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 308898 -2934 309454
rect -2378 308898 19826 309454
rect 20382 308898 55826 309454
rect 56382 308898 91826 309454
rect 92382 308898 127826 309454
rect 128382 308898 163826 309454
rect 164382 308898 199826 309454
rect 200382 308898 235826 309454
rect 236382 308898 271826 309454
rect 272382 308898 307826 309454
rect 308382 308898 343826 309454
rect 344382 308898 379826 309454
rect 380382 308898 415826 309454
rect 416382 308898 451826 309454
rect 452382 308898 487826 309454
rect 488382 308898 523826 309454
rect 524382 308898 559826 309454
rect 560382 308898 586302 309454
rect 586858 308898 586890 309454
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302058 -7734 302614
rect -7178 302058 12986 302614
rect 13542 302058 48986 302614
rect 49542 302058 84986 302614
rect 85542 302058 120986 302614
rect 121542 302058 156986 302614
rect 157542 302058 192986 302614
rect 193542 302058 228986 302614
rect 229542 302058 264986 302614
rect 265542 302058 300986 302614
rect 301542 302058 336986 302614
rect 337542 302058 372986 302614
rect 373542 302058 408986 302614
rect 409542 302058 444986 302614
rect 445542 302058 480986 302614
rect 481542 302058 516986 302614
rect 517542 302058 552986 302614
rect 553542 302058 591102 302614
rect 591658 302058 592650 302614
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298338 -5814 298894
rect -5258 298338 9266 298894
rect 9822 298338 45266 298894
rect 45822 298338 81266 298894
rect 81822 298338 117266 298894
rect 117822 298338 153266 298894
rect 153822 298338 189266 298894
rect 189822 298338 225266 298894
rect 225822 298338 261266 298894
rect 261822 298338 297266 298894
rect 297822 298338 333266 298894
rect 333822 298338 369266 298894
rect 369822 298338 405266 298894
rect 405822 298338 441266 298894
rect 441822 298338 477266 298894
rect 477822 298338 513266 298894
rect 513822 298338 549266 298894
rect 549822 298338 589182 298894
rect 589738 298338 590730 298894
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294618 -3894 295174
rect -3338 294618 5546 295174
rect 6102 294618 41546 295174
rect 42102 294618 77546 295174
rect 78102 294618 113546 295174
rect 114102 294618 149546 295174
rect 150102 294618 185546 295174
rect 186102 294618 221546 295174
rect 222102 294618 257546 295174
rect 258102 294618 293546 295174
rect 294102 294618 329546 295174
rect 330102 294618 365546 295174
rect 366102 294618 401546 295174
rect 402102 294618 437546 295174
rect 438102 294618 473546 295174
rect 474102 294618 509546 295174
rect 510102 294618 545546 295174
rect 546102 294618 581546 295174
rect 582102 294618 587262 295174
rect 587818 294618 588810 295174
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 290898 -1974 291454
rect -1418 290898 1826 291454
rect 2382 290898 37826 291454
rect 38382 290898 73826 291454
rect 74382 290898 109826 291454
rect 110382 290898 145826 291454
rect 146382 290898 181826 291454
rect 182382 290898 217826 291454
rect 218382 290898 253826 291454
rect 254382 290898 289826 291454
rect 290382 290898 325826 291454
rect 326382 290898 361826 291454
rect 362382 290898 397826 291454
rect 398382 290898 433826 291454
rect 434382 290898 469826 291454
rect 470382 290898 505826 291454
rect 506382 290898 541826 291454
rect 542382 290898 577826 291454
rect 578382 290898 585342 291454
rect 585898 290898 586890 291454
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284058 -8694 284614
rect -8138 284058 30986 284614
rect 31542 284058 66986 284614
rect 67542 284058 102986 284614
rect 103542 284058 138986 284614
rect 139542 284058 174986 284614
rect 175542 284058 210986 284614
rect 211542 284058 246986 284614
rect 247542 284058 282986 284614
rect 283542 284058 318986 284614
rect 319542 284058 354986 284614
rect 355542 284058 390986 284614
rect 391542 284058 426986 284614
rect 427542 284058 462986 284614
rect 463542 284058 498986 284614
rect 499542 284058 534986 284614
rect 535542 284058 570986 284614
rect 571542 284058 592062 284614
rect 592618 284058 592650 284614
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280338 -6774 280894
rect -6218 280338 27266 280894
rect 27822 280338 63266 280894
rect 63822 280338 99266 280894
rect 99822 280338 135266 280894
rect 135822 280338 171266 280894
rect 171822 280338 207266 280894
rect 207822 280338 243266 280894
rect 243822 280338 279266 280894
rect 279822 280338 315266 280894
rect 315822 280338 351266 280894
rect 351822 280338 387266 280894
rect 387822 280338 423266 280894
rect 423822 280338 459266 280894
rect 459822 280338 495266 280894
rect 495822 280338 531266 280894
rect 531822 280338 567266 280894
rect 567822 280338 590142 280894
rect 590698 280338 590730 280894
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276618 -4854 277174
rect -4298 276618 23546 277174
rect 24102 276618 59546 277174
rect 60102 276618 95546 277174
rect 96102 276618 131546 277174
rect 132102 276618 167546 277174
rect 168102 276618 203546 277174
rect 204102 276618 239546 277174
rect 240102 276618 275546 277174
rect 276102 276618 311546 277174
rect 312102 276618 347546 277174
rect 348102 276618 383546 277174
rect 384102 276618 419546 277174
rect 420102 276618 455546 277174
rect 456102 276618 491546 277174
rect 492102 276618 527546 277174
rect 528102 276618 563546 277174
rect 564102 276618 588222 277174
rect 588778 276618 588810 277174
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 272898 -2934 273454
rect -2378 272898 19826 273454
rect 20382 272898 55826 273454
rect 56382 272898 91826 273454
rect 92382 272898 127826 273454
rect 128382 272898 163826 273454
rect 164382 272898 199826 273454
rect 200382 272898 235826 273454
rect 236382 272898 271826 273454
rect 272382 272898 307826 273454
rect 308382 272898 343826 273454
rect 344382 272898 379826 273454
rect 380382 272898 415826 273454
rect 416382 272898 451826 273454
rect 452382 272898 487826 273454
rect 488382 272898 523826 273454
rect 524382 272898 559826 273454
rect 560382 272898 586302 273454
rect 586858 272898 586890 273454
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266058 -7734 266614
rect -7178 266058 12986 266614
rect 13542 266058 48986 266614
rect 49542 266058 84986 266614
rect 85542 266058 120986 266614
rect 121542 266058 156986 266614
rect 157542 266058 192986 266614
rect 193542 266058 228986 266614
rect 229542 266058 264986 266614
rect 265542 266058 300986 266614
rect 301542 266058 336986 266614
rect 337542 266058 372986 266614
rect 373542 266058 408986 266614
rect 409542 266058 444986 266614
rect 445542 266058 480986 266614
rect 481542 266058 516986 266614
rect 517542 266058 552986 266614
rect 553542 266058 591102 266614
rect 591658 266058 592650 266614
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262338 -5814 262894
rect -5258 262338 9266 262894
rect 9822 262338 45266 262894
rect 45822 262338 81266 262894
rect 81822 262338 117266 262894
rect 117822 262338 153266 262894
rect 153822 262338 189266 262894
rect 189822 262338 225266 262894
rect 225822 262338 261266 262894
rect 261822 262338 297266 262894
rect 297822 262338 333266 262894
rect 333822 262338 369266 262894
rect 369822 262338 405266 262894
rect 405822 262338 441266 262894
rect 441822 262338 477266 262894
rect 477822 262338 513266 262894
rect 513822 262338 549266 262894
rect 549822 262338 589182 262894
rect 589738 262338 590730 262894
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258618 -3894 259174
rect -3338 258618 5546 259174
rect 6102 258618 41546 259174
rect 42102 258618 77546 259174
rect 78102 258618 113546 259174
rect 114102 258618 149546 259174
rect 150102 258618 185546 259174
rect 186102 258618 221546 259174
rect 222102 258618 257546 259174
rect 258102 258618 293546 259174
rect 294102 258618 329546 259174
rect 330102 258618 365546 259174
rect 366102 258618 401546 259174
rect 402102 258618 437546 259174
rect 438102 258618 473546 259174
rect 474102 258618 509546 259174
rect 510102 258618 545546 259174
rect 546102 258618 581546 259174
rect 582102 258618 587262 259174
rect 587818 258618 588810 259174
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 254898 -1974 255454
rect -1418 254898 1826 255454
rect 2382 254898 37826 255454
rect 38382 254898 73826 255454
rect 74382 254898 109826 255454
rect 110382 254898 145826 255454
rect 146382 254898 181826 255454
rect 182382 254898 217826 255454
rect 218382 254898 253826 255454
rect 254382 254898 289826 255454
rect 290382 254898 325826 255454
rect 326382 254898 361826 255454
rect 362382 254898 397826 255454
rect 398382 254898 433826 255454
rect 434382 254898 469826 255454
rect 470382 254898 505826 255454
rect 506382 254898 541826 255454
rect 542382 254898 577826 255454
rect 578382 254898 585342 255454
rect 585898 254898 586890 255454
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248058 -8694 248614
rect -8138 248058 30986 248614
rect 31542 248058 66986 248614
rect 67542 248058 102986 248614
rect 103542 248058 138986 248614
rect 139542 248058 174986 248614
rect 175542 248058 210986 248614
rect 211542 248058 246986 248614
rect 247542 248058 282986 248614
rect 283542 248058 318986 248614
rect 319542 248058 354986 248614
rect 355542 248058 390986 248614
rect 391542 248058 426986 248614
rect 427542 248058 462986 248614
rect 463542 248058 498986 248614
rect 499542 248058 534986 248614
rect 535542 248058 570986 248614
rect 571542 248058 592062 248614
rect 592618 248058 592650 248614
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244338 -6774 244894
rect -6218 244338 27266 244894
rect 27822 244338 63266 244894
rect 63822 244338 99266 244894
rect 99822 244338 135266 244894
rect 135822 244338 171266 244894
rect 171822 244338 207266 244894
rect 207822 244338 243266 244894
rect 243822 244338 279266 244894
rect 279822 244338 315266 244894
rect 315822 244338 351266 244894
rect 351822 244338 387266 244894
rect 387822 244338 423266 244894
rect 423822 244338 459266 244894
rect 459822 244338 495266 244894
rect 495822 244338 531266 244894
rect 531822 244338 567266 244894
rect 567822 244338 590142 244894
rect 590698 244338 590730 244894
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240618 -4854 241174
rect -4298 240618 23546 241174
rect 24102 240618 59546 241174
rect 60102 240618 95546 241174
rect 96102 240618 131546 241174
rect 132102 240618 167546 241174
rect 168102 240618 203546 241174
rect 204102 240618 239546 241174
rect 240102 240618 275546 241174
rect 276102 240618 311546 241174
rect 312102 240618 347546 241174
rect 348102 240618 383546 241174
rect 384102 240618 419546 241174
rect 420102 240618 455546 241174
rect 456102 240618 491546 241174
rect 492102 240618 527546 241174
rect 528102 240618 563546 241174
rect 564102 240618 588222 241174
rect 588778 240618 588810 241174
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 236898 -2934 237454
rect -2378 236898 19826 237454
rect 20382 236898 55826 237454
rect 56382 236898 91826 237454
rect 92382 236898 127826 237454
rect 128382 236898 163826 237454
rect 164382 236898 199826 237454
rect 200382 236898 235826 237454
rect 236382 236898 271826 237454
rect 272382 236898 307826 237454
rect 308382 236898 343826 237454
rect 344382 236898 379826 237454
rect 380382 236898 415826 237454
rect 416382 236898 451826 237454
rect 452382 236898 487826 237454
rect 488382 236898 523826 237454
rect 524382 236898 559826 237454
rect 560382 236898 586302 237454
rect 586858 236898 586890 237454
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230058 -7734 230614
rect -7178 230058 12986 230614
rect 13542 230058 48986 230614
rect 49542 230058 84986 230614
rect 85542 230058 120986 230614
rect 121542 230058 156986 230614
rect 157542 230058 192986 230614
rect 193542 230058 228986 230614
rect 229542 230058 264986 230614
rect 265542 230058 300986 230614
rect 301542 230058 336986 230614
rect 337542 230058 372986 230614
rect 373542 230058 408986 230614
rect 409542 230058 444986 230614
rect 445542 230058 480986 230614
rect 481542 230058 516986 230614
rect 517542 230058 552986 230614
rect 553542 230058 591102 230614
rect 591658 230058 592650 230614
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226338 -5814 226894
rect -5258 226338 9266 226894
rect 9822 226338 45266 226894
rect 45822 226338 81266 226894
rect 81822 226338 117266 226894
rect 117822 226338 153266 226894
rect 153822 226338 189266 226894
rect 189822 226338 225266 226894
rect 225822 226338 261266 226894
rect 261822 226338 297266 226894
rect 297822 226338 333266 226894
rect 333822 226338 369266 226894
rect 369822 226338 405266 226894
rect 405822 226338 441266 226894
rect 441822 226338 477266 226894
rect 477822 226338 513266 226894
rect 513822 226338 549266 226894
rect 549822 226338 589182 226894
rect 589738 226338 590730 226894
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222618 -3894 223174
rect -3338 222618 5546 223174
rect 6102 222618 41546 223174
rect 42102 222618 77546 223174
rect 78102 222618 113546 223174
rect 114102 222618 149546 223174
rect 150102 222618 185546 223174
rect 186102 222618 221546 223174
rect 222102 222618 257546 223174
rect 258102 222618 293546 223174
rect 294102 222618 329546 223174
rect 330102 222618 365546 223174
rect 366102 222618 401546 223174
rect 402102 222618 437546 223174
rect 438102 222618 473546 223174
rect 474102 222618 509546 223174
rect 510102 222618 545546 223174
rect 546102 222618 581546 223174
rect 582102 222618 587262 223174
rect 587818 222618 588810 223174
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 218898 -1974 219454
rect -1418 218898 1826 219454
rect 2382 218898 37826 219454
rect 38382 218898 73826 219454
rect 74382 218898 109826 219454
rect 110382 218898 145826 219454
rect 146382 218898 181826 219454
rect 182382 218898 217826 219454
rect 218382 218898 253826 219454
rect 254382 218898 289826 219454
rect 290382 218898 325826 219454
rect 326382 218898 361826 219454
rect 362382 218898 397826 219454
rect 398382 218898 433826 219454
rect 434382 218898 469826 219454
rect 470382 218898 505826 219454
rect 506382 218898 541826 219454
rect 542382 218898 577826 219454
rect 578382 218898 585342 219454
rect 585898 218898 586890 219454
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212058 -8694 212614
rect -8138 212058 30986 212614
rect 31542 212058 66986 212614
rect 67542 212058 102986 212614
rect 103542 212058 138986 212614
rect 139542 212058 174986 212614
rect 175542 212058 210986 212614
rect 211542 212058 246986 212614
rect 247542 212058 282986 212614
rect 283542 212058 318986 212614
rect 319542 212058 354986 212614
rect 355542 212058 390986 212614
rect 391542 212058 426986 212614
rect 427542 212058 462986 212614
rect 463542 212058 498986 212614
rect 499542 212058 534986 212614
rect 535542 212058 570986 212614
rect 571542 212058 592062 212614
rect 592618 212058 592650 212614
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208338 -6774 208894
rect -6218 208338 27266 208894
rect 27822 208338 63266 208894
rect 63822 208338 99266 208894
rect 99822 208338 135266 208894
rect 135822 208338 171266 208894
rect 171822 208338 207266 208894
rect 207822 208338 243266 208894
rect 243822 208338 279266 208894
rect 279822 208338 315266 208894
rect 315822 208338 351266 208894
rect 351822 208338 387266 208894
rect 387822 208338 423266 208894
rect 423822 208338 459266 208894
rect 459822 208338 495266 208894
rect 495822 208338 531266 208894
rect 531822 208338 567266 208894
rect 567822 208338 590142 208894
rect 590698 208338 590730 208894
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204618 -4854 205174
rect -4298 204618 23546 205174
rect 24102 204618 59546 205174
rect 60102 204618 95546 205174
rect 96102 204618 131546 205174
rect 132102 204618 167546 205174
rect 168102 204618 203546 205174
rect 204102 204618 239546 205174
rect 240102 204618 275546 205174
rect 276102 204618 311546 205174
rect 312102 204618 347546 205174
rect 348102 204618 383546 205174
rect 384102 204618 419546 205174
rect 420102 204618 455546 205174
rect 456102 204618 491546 205174
rect 492102 204618 527546 205174
rect 528102 204618 563546 205174
rect 564102 204618 588222 205174
rect 588778 204618 588810 205174
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 200898 -2934 201454
rect -2378 200898 19826 201454
rect 20382 200898 55826 201454
rect 56382 200898 91826 201454
rect 92382 200898 127826 201454
rect 128382 200898 163826 201454
rect 164382 200898 199826 201454
rect 200382 200898 235826 201454
rect 236382 200898 271826 201454
rect 272382 200898 307826 201454
rect 308382 200898 343826 201454
rect 344382 200898 379826 201454
rect 380382 200898 415826 201454
rect 416382 200898 451826 201454
rect 452382 200898 487826 201454
rect 488382 200898 523826 201454
rect 524382 200898 559826 201454
rect 560382 200898 586302 201454
rect 586858 200898 586890 201454
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194058 -7734 194614
rect -7178 194058 12986 194614
rect 13542 194058 48986 194614
rect 49542 194058 84986 194614
rect 85542 194058 120986 194614
rect 121542 194058 156986 194614
rect 157542 194058 192986 194614
rect 193542 194058 228986 194614
rect 229542 194058 264986 194614
rect 265542 194058 300986 194614
rect 301542 194058 336986 194614
rect 337542 194058 372986 194614
rect 373542 194058 408986 194614
rect 409542 194058 444986 194614
rect 445542 194058 480986 194614
rect 481542 194058 516986 194614
rect 517542 194058 552986 194614
rect 553542 194058 591102 194614
rect 591658 194058 592650 194614
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190338 -5814 190894
rect -5258 190338 9266 190894
rect 9822 190338 45266 190894
rect 45822 190338 81266 190894
rect 81822 190338 117266 190894
rect 117822 190338 153266 190894
rect 153822 190338 189266 190894
rect 189822 190338 225266 190894
rect 225822 190338 261266 190894
rect 261822 190338 297266 190894
rect 297822 190338 333266 190894
rect 333822 190338 369266 190894
rect 369822 190338 405266 190894
rect 405822 190338 441266 190894
rect 441822 190338 477266 190894
rect 477822 190338 513266 190894
rect 513822 190338 549266 190894
rect 549822 190338 589182 190894
rect 589738 190338 590730 190894
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186618 -3894 187174
rect -3338 186618 5546 187174
rect 6102 186618 41546 187174
rect 42102 186618 77546 187174
rect 78102 186618 113546 187174
rect 114102 186618 149546 187174
rect 150102 186618 185546 187174
rect 186102 186618 221546 187174
rect 222102 186618 257546 187174
rect 258102 186618 293546 187174
rect 294102 186618 329546 187174
rect 330102 186618 365546 187174
rect 366102 186618 401546 187174
rect 402102 186618 437546 187174
rect 438102 186618 473546 187174
rect 474102 186618 509546 187174
rect 510102 186618 545546 187174
rect 546102 186618 581546 187174
rect 582102 186618 587262 187174
rect 587818 186618 588810 187174
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 182898 -1974 183454
rect -1418 182898 1826 183454
rect 2382 182898 37826 183454
rect 38382 182898 73826 183454
rect 74382 182898 109826 183454
rect 110382 182898 145826 183454
rect 146382 182898 181826 183454
rect 182382 182898 217826 183454
rect 218382 182898 253826 183454
rect 254382 182898 289826 183454
rect 290382 182898 325826 183454
rect 326382 182898 361826 183454
rect 362382 182898 397826 183454
rect 398382 182898 433826 183454
rect 434382 182898 469826 183454
rect 470382 182898 505826 183454
rect 506382 182898 541826 183454
rect 542382 182898 577826 183454
rect 578382 182898 585342 183454
rect 585898 182898 586890 183454
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176058 -8694 176614
rect -8138 176058 30986 176614
rect 31542 176058 66986 176614
rect 67542 176058 102986 176614
rect 103542 176058 138986 176614
rect 139542 176058 174986 176614
rect 175542 176058 210986 176614
rect 211542 176058 246986 176614
rect 247542 176058 282986 176614
rect 283542 176058 318986 176614
rect 319542 176058 354986 176614
rect 355542 176058 390986 176614
rect 391542 176058 426986 176614
rect 427542 176058 462986 176614
rect 463542 176058 498986 176614
rect 499542 176058 534986 176614
rect 535542 176058 570986 176614
rect 571542 176058 592062 176614
rect 592618 176058 592650 176614
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172338 -6774 172894
rect -6218 172338 27266 172894
rect 27822 172338 63266 172894
rect 63822 172338 99266 172894
rect 99822 172338 135266 172894
rect 135822 172338 171266 172894
rect 171822 172338 207266 172894
rect 207822 172338 243266 172894
rect 243822 172338 279266 172894
rect 279822 172338 315266 172894
rect 315822 172338 351266 172894
rect 351822 172338 387266 172894
rect 387822 172338 423266 172894
rect 423822 172338 459266 172894
rect 459822 172338 495266 172894
rect 495822 172338 531266 172894
rect 531822 172338 567266 172894
rect 567822 172338 590142 172894
rect 590698 172338 590730 172894
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168618 -4854 169174
rect -4298 168618 23546 169174
rect 24102 168618 59546 169174
rect 60102 168618 95546 169174
rect 96102 168618 131546 169174
rect 132102 168618 167546 169174
rect 168102 168618 203546 169174
rect 204102 168618 239546 169174
rect 240102 168618 275546 169174
rect 276102 168618 311546 169174
rect 312102 168618 347546 169174
rect 348102 168618 383546 169174
rect 384102 168618 419546 169174
rect 420102 168618 455546 169174
rect 456102 168618 491546 169174
rect 492102 168618 527546 169174
rect 528102 168618 563546 169174
rect 564102 168618 588222 169174
rect 588778 168618 588810 169174
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 164898 -2934 165454
rect -2378 164898 19826 165454
rect 20382 164898 55826 165454
rect 56382 164898 91826 165454
rect 92382 164898 127826 165454
rect 128382 164898 163826 165454
rect 164382 164898 199826 165454
rect 200382 164898 235826 165454
rect 236382 164898 271826 165454
rect 272382 164898 307826 165454
rect 308382 164898 343826 165454
rect 344382 164898 379826 165454
rect 380382 164898 415826 165454
rect 416382 164898 451826 165454
rect 452382 164898 487826 165454
rect 488382 164898 523826 165454
rect 524382 164898 559826 165454
rect 560382 164898 586302 165454
rect 586858 164898 586890 165454
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158058 -7734 158614
rect -7178 158058 12986 158614
rect 13542 158058 48986 158614
rect 49542 158058 84986 158614
rect 85542 158058 120986 158614
rect 121542 158058 156986 158614
rect 157542 158058 192986 158614
rect 193542 158058 228986 158614
rect 229542 158058 264986 158614
rect 265542 158058 300986 158614
rect 301542 158058 336986 158614
rect 337542 158058 372986 158614
rect 373542 158058 408986 158614
rect 409542 158058 444986 158614
rect 445542 158058 480986 158614
rect 481542 158058 516986 158614
rect 517542 158058 552986 158614
rect 553542 158058 591102 158614
rect 591658 158058 592650 158614
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154338 -5814 154894
rect -5258 154338 9266 154894
rect 9822 154338 45266 154894
rect 45822 154338 81266 154894
rect 81822 154338 117266 154894
rect 117822 154338 153266 154894
rect 153822 154338 189266 154894
rect 189822 154338 225266 154894
rect 225822 154338 261266 154894
rect 261822 154338 297266 154894
rect 297822 154338 333266 154894
rect 333822 154338 369266 154894
rect 369822 154338 405266 154894
rect 405822 154338 441266 154894
rect 441822 154338 477266 154894
rect 477822 154338 513266 154894
rect 513822 154338 549266 154894
rect 549822 154338 589182 154894
rect 589738 154338 590730 154894
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150618 -3894 151174
rect -3338 150618 5546 151174
rect 6102 150618 41546 151174
rect 42102 150618 77546 151174
rect 78102 150618 113546 151174
rect 114102 150618 149546 151174
rect 150102 150618 185546 151174
rect 186102 150618 221546 151174
rect 222102 150618 257546 151174
rect 258102 150618 293546 151174
rect 294102 150618 329546 151174
rect 330102 150618 365546 151174
rect 366102 150618 401546 151174
rect 402102 150618 437546 151174
rect 438102 150618 473546 151174
rect 474102 150618 509546 151174
rect 510102 150618 545546 151174
rect 546102 150618 581546 151174
rect 582102 150618 587262 151174
rect 587818 150618 588810 151174
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 146898 -1974 147454
rect -1418 146898 1826 147454
rect 2382 146898 37826 147454
rect 38382 146898 73826 147454
rect 74382 146898 109826 147454
rect 110382 146898 145826 147454
rect 146382 146898 181826 147454
rect 182382 146898 217826 147454
rect 218382 146898 253826 147454
rect 254382 146898 289826 147454
rect 290382 146898 325826 147454
rect 326382 146898 361826 147454
rect 362382 146898 397826 147454
rect 398382 146898 433826 147454
rect 434382 146898 469826 147454
rect 470382 146898 505826 147454
rect 506382 146898 541826 147454
rect 542382 146898 577826 147454
rect 578382 146898 585342 147454
rect 585898 146898 586890 147454
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140058 -8694 140614
rect -8138 140058 30986 140614
rect 31542 140058 66986 140614
rect 67542 140058 102986 140614
rect 103542 140058 138986 140614
rect 139542 140058 174986 140614
rect 175542 140058 210986 140614
rect 211542 140058 246986 140614
rect 247542 140058 282986 140614
rect 283542 140058 318986 140614
rect 319542 140058 354986 140614
rect 355542 140058 390986 140614
rect 391542 140058 426986 140614
rect 427542 140058 462986 140614
rect 463542 140058 498986 140614
rect 499542 140058 534986 140614
rect 535542 140058 570986 140614
rect 571542 140058 592062 140614
rect 592618 140058 592650 140614
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136338 -6774 136894
rect -6218 136338 27266 136894
rect 27822 136338 63266 136894
rect 63822 136338 99266 136894
rect 99822 136338 135266 136894
rect 135822 136338 171266 136894
rect 171822 136338 207266 136894
rect 207822 136338 243266 136894
rect 243822 136338 279266 136894
rect 279822 136338 315266 136894
rect 315822 136338 351266 136894
rect 351822 136338 387266 136894
rect 387822 136338 423266 136894
rect 423822 136338 459266 136894
rect 459822 136338 495266 136894
rect 495822 136338 531266 136894
rect 531822 136338 567266 136894
rect 567822 136338 590142 136894
rect 590698 136338 590730 136894
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132618 -4854 133174
rect -4298 132618 23546 133174
rect 24102 132618 59546 133174
rect 60102 132618 95546 133174
rect 96102 132618 131546 133174
rect 132102 132618 167546 133174
rect 168102 132618 203546 133174
rect 204102 132618 239546 133174
rect 240102 132618 275546 133174
rect 276102 132618 311546 133174
rect 312102 132618 347546 133174
rect 348102 132618 383546 133174
rect 384102 132618 419546 133174
rect 420102 132618 455546 133174
rect 456102 132618 491546 133174
rect 492102 132618 527546 133174
rect 528102 132618 563546 133174
rect 564102 132618 588222 133174
rect 588778 132618 588810 133174
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 128898 -2934 129454
rect -2378 128898 19826 129454
rect 20382 128898 55826 129454
rect 56382 128898 91826 129454
rect 92382 128898 127826 129454
rect 128382 128898 163826 129454
rect 164382 128898 199826 129454
rect 200382 128898 235826 129454
rect 236382 128898 271826 129454
rect 272382 128898 307826 129454
rect 308382 128898 343826 129454
rect 344382 128898 379826 129454
rect 380382 128898 415826 129454
rect 416382 128898 451826 129454
rect 452382 128898 487826 129454
rect 488382 128898 523826 129454
rect 524382 128898 559826 129454
rect 560382 128898 586302 129454
rect 586858 128898 586890 129454
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122058 -7734 122614
rect -7178 122058 12986 122614
rect 13542 122058 48986 122614
rect 49542 122058 84986 122614
rect 85542 122058 120986 122614
rect 121542 122058 156986 122614
rect 157542 122058 192986 122614
rect 193542 122058 228986 122614
rect 229542 122058 264986 122614
rect 265542 122058 300986 122614
rect 301542 122058 336986 122614
rect 337542 122058 372986 122614
rect 373542 122058 408986 122614
rect 409542 122058 444986 122614
rect 445542 122058 480986 122614
rect 481542 122058 516986 122614
rect 517542 122058 552986 122614
rect 553542 122058 591102 122614
rect 591658 122058 592650 122614
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118338 -5814 118894
rect -5258 118338 9266 118894
rect 9822 118338 45266 118894
rect 45822 118338 81266 118894
rect 81822 118338 117266 118894
rect 117822 118338 153266 118894
rect 153822 118338 189266 118894
rect 189822 118338 225266 118894
rect 225822 118338 261266 118894
rect 261822 118338 297266 118894
rect 297822 118338 333266 118894
rect 333822 118338 369266 118894
rect 369822 118338 405266 118894
rect 405822 118338 441266 118894
rect 441822 118338 477266 118894
rect 477822 118338 513266 118894
rect 513822 118338 549266 118894
rect 549822 118338 589182 118894
rect 589738 118338 590730 118894
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114618 -3894 115174
rect -3338 114618 5546 115174
rect 6102 114618 41546 115174
rect 42102 114618 77546 115174
rect 78102 114618 113546 115174
rect 114102 114618 149546 115174
rect 150102 114618 185546 115174
rect 186102 114618 221546 115174
rect 222102 114618 257546 115174
rect 258102 114618 293546 115174
rect 294102 114618 329546 115174
rect 330102 114618 365546 115174
rect 366102 114618 401546 115174
rect 402102 114618 437546 115174
rect 438102 114618 473546 115174
rect 474102 114618 509546 115174
rect 510102 114618 545546 115174
rect 546102 114618 581546 115174
rect 582102 114618 587262 115174
rect 587818 114618 588810 115174
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 110898 -1974 111454
rect -1418 110898 1826 111454
rect 2382 110898 37826 111454
rect 38382 110898 73826 111454
rect 74382 110898 109826 111454
rect 110382 110898 145826 111454
rect 146382 110898 181826 111454
rect 182382 110898 217826 111454
rect 218382 110898 253826 111454
rect 254382 110898 289826 111454
rect 290382 110898 325826 111454
rect 326382 110898 361826 111454
rect 362382 110898 397826 111454
rect 398382 110898 433826 111454
rect 434382 110898 469826 111454
rect 470382 110898 505826 111454
rect 506382 110898 541826 111454
rect 542382 110898 577826 111454
rect 578382 110898 585342 111454
rect 585898 110898 586890 111454
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104058 -8694 104614
rect -8138 104058 30986 104614
rect 31542 104058 66986 104614
rect 67542 104058 102986 104614
rect 103542 104058 138986 104614
rect 139542 104058 174986 104614
rect 175542 104058 210986 104614
rect 211542 104058 246986 104614
rect 247542 104058 282986 104614
rect 283542 104058 318986 104614
rect 319542 104058 354986 104614
rect 355542 104058 390986 104614
rect 391542 104058 426986 104614
rect 427542 104058 462986 104614
rect 463542 104058 498986 104614
rect 499542 104058 534986 104614
rect 535542 104058 570986 104614
rect 571542 104058 592062 104614
rect 592618 104058 592650 104614
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100338 -6774 100894
rect -6218 100338 27266 100894
rect 27822 100338 63266 100894
rect 63822 100338 99266 100894
rect 99822 100338 135266 100894
rect 135822 100338 171266 100894
rect 171822 100338 207266 100894
rect 207822 100338 243266 100894
rect 243822 100338 279266 100894
rect 279822 100338 315266 100894
rect 315822 100338 351266 100894
rect 351822 100338 387266 100894
rect 387822 100338 423266 100894
rect 423822 100338 459266 100894
rect 459822 100338 495266 100894
rect 495822 100338 531266 100894
rect 531822 100338 567266 100894
rect 567822 100338 590142 100894
rect 590698 100338 590730 100894
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96618 -4854 97174
rect -4298 96618 23546 97174
rect 24102 96618 59546 97174
rect 60102 96618 95546 97174
rect 96102 96618 131546 97174
rect 132102 96618 167546 97174
rect 168102 96618 203546 97174
rect 204102 96618 239546 97174
rect 240102 96618 275546 97174
rect 276102 96618 311546 97174
rect 312102 96618 347546 97174
rect 348102 96618 383546 97174
rect 384102 96618 419546 97174
rect 420102 96618 455546 97174
rect 456102 96618 491546 97174
rect 492102 96618 527546 97174
rect 528102 96618 563546 97174
rect 564102 96618 588222 97174
rect 588778 96618 588810 97174
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 92898 -2934 93454
rect -2378 92898 19826 93454
rect 20382 92898 55826 93454
rect 56382 92898 91826 93454
rect 92382 92898 127826 93454
rect 128382 92898 163826 93454
rect 164382 92898 199826 93454
rect 200382 92898 235826 93454
rect 236382 92898 271826 93454
rect 272382 92898 307826 93454
rect 308382 92898 343826 93454
rect 344382 92898 379826 93454
rect 380382 92898 415826 93454
rect 416382 92898 451826 93454
rect 452382 92898 487826 93454
rect 488382 92898 523826 93454
rect 524382 92898 559826 93454
rect 560382 92898 586302 93454
rect 586858 92898 586890 93454
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86058 -7734 86614
rect -7178 86058 12986 86614
rect 13542 86058 48986 86614
rect 49542 86058 84986 86614
rect 85542 86058 120986 86614
rect 121542 86058 156986 86614
rect 157542 86058 192986 86614
rect 193542 86058 228986 86614
rect 229542 86058 264986 86614
rect 265542 86058 300986 86614
rect 301542 86058 336986 86614
rect 337542 86058 372986 86614
rect 373542 86058 408986 86614
rect 409542 86058 444986 86614
rect 445542 86058 480986 86614
rect 481542 86058 516986 86614
rect 517542 86058 552986 86614
rect 553542 86058 591102 86614
rect 591658 86058 592650 86614
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82338 -5814 82894
rect -5258 82338 9266 82894
rect 9822 82338 45266 82894
rect 45822 82338 81266 82894
rect 81822 82338 117266 82894
rect 117822 82338 153266 82894
rect 153822 82338 189266 82894
rect 189822 82338 225266 82894
rect 225822 82338 261266 82894
rect 261822 82338 297266 82894
rect 297822 82338 333266 82894
rect 333822 82338 369266 82894
rect 369822 82338 405266 82894
rect 405822 82338 441266 82894
rect 441822 82338 477266 82894
rect 477822 82338 513266 82894
rect 513822 82338 549266 82894
rect 549822 82338 589182 82894
rect 589738 82338 590730 82894
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78618 -3894 79174
rect -3338 78618 5546 79174
rect 6102 78618 41546 79174
rect 42102 78618 77546 79174
rect 78102 78618 113546 79174
rect 114102 78618 149546 79174
rect 150102 78618 185546 79174
rect 186102 78618 221546 79174
rect 222102 78618 257546 79174
rect 258102 78618 293546 79174
rect 294102 78618 329546 79174
rect 330102 78618 365546 79174
rect 366102 78618 401546 79174
rect 402102 78618 437546 79174
rect 438102 78618 473546 79174
rect 474102 78618 509546 79174
rect 510102 78618 545546 79174
rect 546102 78618 581546 79174
rect 582102 78618 587262 79174
rect 587818 78618 588810 79174
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 74898 -1974 75454
rect -1418 74898 1826 75454
rect 2382 74898 37826 75454
rect 38382 74898 73826 75454
rect 74382 74898 109826 75454
rect 110382 74898 145826 75454
rect 146382 74898 181826 75454
rect 182382 74898 217826 75454
rect 218382 74898 253826 75454
rect 254382 74898 289826 75454
rect 290382 74898 325826 75454
rect 326382 74898 361826 75454
rect 362382 74898 397826 75454
rect 398382 74898 433826 75454
rect 434382 74898 469826 75454
rect 470382 74898 505826 75454
rect 506382 74898 541826 75454
rect 542382 74898 577826 75454
rect 578382 74898 585342 75454
rect 585898 74898 586890 75454
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68058 -8694 68614
rect -8138 68058 30986 68614
rect 31542 68058 66986 68614
rect 67542 68058 102986 68614
rect 103542 68058 138986 68614
rect 139542 68058 174986 68614
rect 175542 68058 210986 68614
rect 211542 68058 246986 68614
rect 247542 68058 282986 68614
rect 283542 68058 318986 68614
rect 319542 68058 354986 68614
rect 355542 68058 390986 68614
rect 391542 68058 426986 68614
rect 427542 68058 462986 68614
rect 463542 68058 498986 68614
rect 499542 68058 534986 68614
rect 535542 68058 570986 68614
rect 571542 68058 592062 68614
rect 592618 68058 592650 68614
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64338 -6774 64894
rect -6218 64338 27266 64894
rect 27822 64338 63266 64894
rect 63822 64338 99266 64894
rect 99822 64338 135266 64894
rect 135822 64338 171266 64894
rect 171822 64338 207266 64894
rect 207822 64338 243266 64894
rect 243822 64338 279266 64894
rect 279822 64338 315266 64894
rect 315822 64338 351266 64894
rect 351822 64338 387266 64894
rect 387822 64338 423266 64894
rect 423822 64338 459266 64894
rect 459822 64338 495266 64894
rect 495822 64338 531266 64894
rect 531822 64338 567266 64894
rect 567822 64338 590142 64894
rect 590698 64338 590730 64894
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60618 -4854 61174
rect -4298 60618 23546 61174
rect 24102 60618 59546 61174
rect 60102 60618 95546 61174
rect 96102 60618 131546 61174
rect 132102 60618 167546 61174
rect 168102 60618 203546 61174
rect 204102 60618 239546 61174
rect 240102 60618 275546 61174
rect 276102 60618 311546 61174
rect 312102 60618 347546 61174
rect 348102 60618 383546 61174
rect 384102 60618 419546 61174
rect 420102 60618 455546 61174
rect 456102 60618 491546 61174
rect 492102 60618 527546 61174
rect 528102 60618 563546 61174
rect 564102 60618 588222 61174
rect 588778 60618 588810 61174
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 56898 -2934 57454
rect -2378 56898 19826 57454
rect 20382 56898 55826 57454
rect 56382 56898 91826 57454
rect 92382 56898 127826 57454
rect 128382 56898 163826 57454
rect 164382 56898 199826 57454
rect 200382 56898 235826 57454
rect 236382 56898 271826 57454
rect 272382 56898 307826 57454
rect 308382 56898 343826 57454
rect 344382 56898 379826 57454
rect 380382 56898 415826 57454
rect 416382 56898 451826 57454
rect 452382 56898 487826 57454
rect 488382 56898 523826 57454
rect 524382 56898 559826 57454
rect 560382 56898 586302 57454
rect 586858 56898 586890 57454
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50058 -7734 50614
rect -7178 50058 12986 50614
rect 13542 50058 48986 50614
rect 49542 50058 84986 50614
rect 85542 50058 120986 50614
rect 121542 50058 156986 50614
rect 157542 50058 192986 50614
rect 193542 50058 228986 50614
rect 229542 50058 264986 50614
rect 265542 50058 300986 50614
rect 301542 50058 336986 50614
rect 337542 50058 372986 50614
rect 373542 50058 408986 50614
rect 409542 50058 444986 50614
rect 445542 50058 480986 50614
rect 481542 50058 516986 50614
rect 517542 50058 552986 50614
rect 553542 50058 591102 50614
rect 591658 50058 592650 50614
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46338 -5814 46894
rect -5258 46338 9266 46894
rect 9822 46338 45266 46894
rect 45822 46338 81266 46894
rect 81822 46338 117266 46894
rect 117822 46338 153266 46894
rect 153822 46338 189266 46894
rect 189822 46338 225266 46894
rect 225822 46338 261266 46894
rect 261822 46338 297266 46894
rect 297822 46338 333266 46894
rect 333822 46338 369266 46894
rect 369822 46338 405266 46894
rect 405822 46338 441266 46894
rect 441822 46338 477266 46894
rect 477822 46338 513266 46894
rect 513822 46338 549266 46894
rect 549822 46338 589182 46894
rect 589738 46338 590730 46894
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42618 -3894 43174
rect -3338 42618 5546 43174
rect 6102 42618 41546 43174
rect 42102 42618 77546 43174
rect 78102 42618 113546 43174
rect 114102 42618 149546 43174
rect 150102 42618 185546 43174
rect 186102 42618 221546 43174
rect 222102 42618 257546 43174
rect 258102 42618 293546 43174
rect 294102 42618 329546 43174
rect 330102 42618 365546 43174
rect 366102 42618 401546 43174
rect 402102 42618 437546 43174
rect 438102 42618 473546 43174
rect 474102 42618 509546 43174
rect 510102 42618 545546 43174
rect 546102 42618 581546 43174
rect 582102 42618 587262 43174
rect 587818 42618 588810 43174
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 38898 -1974 39454
rect -1418 38898 1826 39454
rect 2382 38898 37826 39454
rect 38382 38898 73826 39454
rect 74382 38898 109826 39454
rect 110382 38898 145826 39454
rect 146382 38898 181826 39454
rect 182382 38898 217826 39454
rect 218382 38898 253826 39454
rect 254382 38898 289826 39454
rect 290382 38898 325826 39454
rect 326382 38898 361826 39454
rect 362382 38898 397826 39454
rect 398382 38898 433826 39454
rect 434382 38898 469826 39454
rect 470382 38898 505826 39454
rect 506382 38898 541826 39454
rect 542382 38898 577826 39454
rect 578382 38898 585342 39454
rect 585898 38898 586890 39454
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32058 -8694 32614
rect -8138 32058 30986 32614
rect 31542 32058 66986 32614
rect 67542 32058 102986 32614
rect 103542 32058 138986 32614
rect 139542 32058 174986 32614
rect 175542 32058 210986 32614
rect 211542 32058 246986 32614
rect 247542 32058 282986 32614
rect 283542 32058 318986 32614
rect 319542 32058 354986 32614
rect 355542 32058 390986 32614
rect 391542 32058 426986 32614
rect 427542 32058 462986 32614
rect 463542 32058 498986 32614
rect 499542 32058 534986 32614
rect 535542 32058 570986 32614
rect 571542 32058 592062 32614
rect 592618 32058 592650 32614
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28338 -6774 28894
rect -6218 28338 27266 28894
rect 27822 28338 63266 28894
rect 63822 28338 99266 28894
rect 99822 28338 135266 28894
rect 135822 28338 171266 28894
rect 171822 28338 207266 28894
rect 207822 28338 243266 28894
rect 243822 28338 279266 28894
rect 279822 28338 315266 28894
rect 315822 28338 351266 28894
rect 351822 28338 387266 28894
rect 387822 28338 423266 28894
rect 423822 28338 459266 28894
rect 459822 28338 495266 28894
rect 495822 28338 531266 28894
rect 531822 28338 567266 28894
rect 567822 28338 590142 28894
rect 590698 28338 590730 28894
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24618 -4854 25174
rect -4298 24618 23546 25174
rect 24102 24618 59546 25174
rect 60102 24618 95546 25174
rect 96102 24618 131546 25174
rect 132102 24618 167546 25174
rect 168102 24618 203546 25174
rect 204102 24618 239546 25174
rect 240102 24618 275546 25174
rect 276102 24618 311546 25174
rect 312102 24618 347546 25174
rect 348102 24618 383546 25174
rect 384102 24618 419546 25174
rect 420102 24618 455546 25174
rect 456102 24618 491546 25174
rect 492102 24618 527546 25174
rect 528102 24618 563546 25174
rect 564102 24618 588222 25174
rect 588778 24618 588810 25174
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 20898 -2934 21454
rect -2378 20898 19826 21454
rect 20382 20898 55826 21454
rect 56382 20898 91826 21454
rect 92382 20898 127826 21454
rect 128382 20898 163826 21454
rect 164382 20898 199826 21454
rect 200382 20898 235826 21454
rect 236382 20898 271826 21454
rect 272382 20898 307826 21454
rect 308382 20898 343826 21454
rect 344382 20898 379826 21454
rect 380382 20898 415826 21454
rect 416382 20898 451826 21454
rect 452382 20898 487826 21454
rect 488382 20898 523826 21454
rect 524382 20898 559826 21454
rect 560382 20898 586302 21454
rect 586858 20898 586890 21454
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14058 -7734 14614
rect -7178 14058 12986 14614
rect 13542 14058 48986 14614
rect 49542 14058 84986 14614
rect 85542 14058 120986 14614
rect 121542 14058 156986 14614
rect 157542 14058 192986 14614
rect 193542 14058 228986 14614
rect 229542 14058 264986 14614
rect 265542 14058 300986 14614
rect 301542 14058 336986 14614
rect 337542 14058 372986 14614
rect 373542 14058 408986 14614
rect 409542 14058 444986 14614
rect 445542 14058 480986 14614
rect 481542 14058 516986 14614
rect 517542 14058 552986 14614
rect 553542 14058 591102 14614
rect 591658 14058 592650 14614
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10338 -5814 10894
rect -5258 10338 9266 10894
rect 9822 10338 45266 10894
rect 45822 10338 81266 10894
rect 81822 10338 117266 10894
rect 117822 10338 153266 10894
rect 153822 10338 189266 10894
rect 189822 10338 225266 10894
rect 225822 10338 261266 10894
rect 261822 10338 297266 10894
rect 297822 10338 333266 10894
rect 333822 10338 369266 10894
rect 369822 10338 405266 10894
rect 405822 10338 441266 10894
rect 441822 10338 477266 10894
rect 477822 10338 513266 10894
rect 513822 10338 549266 10894
rect 549822 10338 589182 10894
rect 589738 10338 590730 10894
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6618 -3894 7174
rect -3338 6618 5546 7174
rect 6102 6618 41546 7174
rect 42102 6618 77546 7174
rect 78102 6618 113546 7174
rect 114102 6618 149546 7174
rect 150102 6618 185546 7174
rect 186102 6618 221546 7174
rect 222102 6618 257546 7174
rect 258102 6618 293546 7174
rect 294102 6618 329546 7174
rect 330102 6618 365546 7174
rect 366102 6618 401546 7174
rect 402102 6618 437546 7174
rect 438102 6618 473546 7174
rect 474102 6618 509546 7174
rect 510102 6618 545546 7174
rect 546102 6618 581546 7174
rect 582102 6618 587262 7174
rect 587818 6618 588810 7174
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 2898 -1974 3454
rect -1418 2898 1826 3454
rect 2382 2898 37826 3454
rect 38382 2898 73826 3454
rect 74382 2898 109826 3454
rect 110382 2898 145826 3454
rect 146382 2898 181826 3454
rect 182382 2898 217826 3454
rect 218382 2898 253826 3454
rect 254382 2898 289826 3454
rect 290382 2898 325826 3454
rect 326382 2898 361826 3454
rect 362382 2898 397826 3454
rect 398382 2898 433826 3454
rect 434382 2898 469826 3454
rect 470382 2898 505826 3454
rect 506382 2898 541826 3454
rect 542382 2898 577826 3454
rect 578382 2898 585342 3454
rect 585898 2898 586890 3454
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -902 -1974 -346
rect -1418 -902 1826 -346
rect 2382 -902 37826 -346
rect 38382 -902 73826 -346
rect 74382 -902 109826 -346
rect 110382 -902 145826 -346
rect 146382 -902 181826 -346
rect 182382 -902 217826 -346
rect 218382 -902 253826 -346
rect 254382 -902 289826 -346
rect 290382 -902 325826 -346
rect 326382 -902 361826 -346
rect 362382 -902 397826 -346
rect 398382 -902 433826 -346
rect 434382 -902 469826 -346
rect 470382 -902 505826 -346
rect 506382 -902 541826 -346
rect 542382 -902 577826 -346
rect 578382 -902 585342 -346
rect 585898 -902 585930 -346
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1862 -2934 -1306
rect -2378 -1862 19826 -1306
rect 20382 -1862 55826 -1306
rect 56382 -1862 91826 -1306
rect 92382 -1862 127826 -1306
rect 128382 -1862 163826 -1306
rect 164382 -1862 199826 -1306
rect 200382 -1862 235826 -1306
rect 236382 -1862 271826 -1306
rect 272382 -1862 307826 -1306
rect 308382 -1862 343826 -1306
rect 344382 -1862 379826 -1306
rect 380382 -1862 415826 -1306
rect 416382 -1862 451826 -1306
rect 452382 -1862 487826 -1306
rect 488382 -1862 523826 -1306
rect 524382 -1862 559826 -1306
rect 560382 -1862 586302 -1306
rect 586858 -1862 586890 -1306
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2822 -3894 -2266
rect -3338 -2822 5546 -2266
rect 6102 -2822 41546 -2266
rect 42102 -2822 77546 -2266
rect 78102 -2822 113546 -2266
rect 114102 -2822 149546 -2266
rect 150102 -2822 185546 -2266
rect 186102 -2822 221546 -2266
rect 222102 -2822 257546 -2266
rect 258102 -2822 293546 -2266
rect 294102 -2822 329546 -2266
rect 330102 -2822 365546 -2266
rect 366102 -2822 401546 -2266
rect 402102 -2822 437546 -2266
rect 438102 -2822 473546 -2266
rect 474102 -2822 509546 -2266
rect 510102 -2822 545546 -2266
rect 546102 -2822 581546 -2266
rect 582102 -2822 587262 -2266
rect 587818 -2822 587850 -2266
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3782 -4854 -3226
rect -4298 -3782 23546 -3226
rect 24102 -3782 59546 -3226
rect 60102 -3782 95546 -3226
rect 96102 -3782 131546 -3226
rect 132102 -3782 167546 -3226
rect 168102 -3782 203546 -3226
rect 204102 -3782 239546 -3226
rect 240102 -3782 275546 -3226
rect 276102 -3782 311546 -3226
rect 312102 -3782 347546 -3226
rect 348102 -3782 383546 -3226
rect 384102 -3782 419546 -3226
rect 420102 -3782 455546 -3226
rect 456102 -3782 491546 -3226
rect 492102 -3782 527546 -3226
rect 528102 -3782 563546 -3226
rect 564102 -3782 588222 -3226
rect 588778 -3782 588810 -3226
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4742 -5814 -4186
rect -5258 -4742 9266 -4186
rect 9822 -4742 45266 -4186
rect 45822 -4742 81266 -4186
rect 81822 -4742 117266 -4186
rect 117822 -4742 153266 -4186
rect 153822 -4742 189266 -4186
rect 189822 -4742 225266 -4186
rect 225822 -4742 261266 -4186
rect 261822 -4742 297266 -4186
rect 297822 -4742 333266 -4186
rect 333822 -4742 369266 -4186
rect 369822 -4742 405266 -4186
rect 405822 -4742 441266 -4186
rect 441822 -4742 477266 -4186
rect 477822 -4742 513266 -4186
rect 513822 -4742 549266 -4186
rect 549822 -4742 589182 -4186
rect 589738 -4742 589770 -4186
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5702 -6774 -5146
rect -6218 -5702 27266 -5146
rect 27822 -5702 63266 -5146
rect 63822 -5702 99266 -5146
rect 99822 -5702 135266 -5146
rect 135822 -5702 171266 -5146
rect 171822 -5702 207266 -5146
rect 207822 -5702 243266 -5146
rect 243822 -5702 279266 -5146
rect 279822 -5702 315266 -5146
rect 315822 -5702 351266 -5146
rect 351822 -5702 387266 -5146
rect 387822 -5702 423266 -5146
rect 423822 -5702 459266 -5146
rect 459822 -5702 495266 -5146
rect 495822 -5702 531266 -5146
rect 531822 -5702 567266 -5146
rect 567822 -5702 590142 -5146
rect 590698 -5702 590730 -5146
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6662 -7734 -6106
rect -7178 -6662 12986 -6106
rect 13542 -6662 48986 -6106
rect 49542 -6662 84986 -6106
rect 85542 -6662 120986 -6106
rect 121542 -6662 156986 -6106
rect 157542 -6662 192986 -6106
rect 193542 -6662 228986 -6106
rect 229542 -6662 264986 -6106
rect 265542 -6662 300986 -6106
rect 301542 -6662 336986 -6106
rect 337542 -6662 372986 -6106
rect 373542 -6662 408986 -6106
rect 409542 -6662 444986 -6106
rect 445542 -6662 480986 -6106
rect 481542 -6662 516986 -6106
rect 517542 -6662 552986 -6106
rect 553542 -6662 591102 -6106
rect 591658 -6662 591690 -6106
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7622 -8694 -7066
rect -8138 -7622 30986 -7066
rect 31542 -7622 66986 -7066
rect 67542 -7622 102986 -7066
rect 103542 -7622 138986 -7066
rect 139542 -7622 174986 -7066
rect 175542 -7622 210986 -7066
rect 211542 -7622 246986 -7066
rect 247542 -7622 282986 -7066
rect 283542 -7622 318986 -7066
rect 319542 -7622 354986 -7066
rect 355542 -7622 390986 -7066
rect 391542 -7622 426986 -7066
rect 427542 -7622 462986 -7066
rect 463542 -7622 498986 -7066
rect 499542 -7622 534986 -7066
rect 535542 -7622 570986 -7066
rect 571542 -7622 592062 -7066
rect 592618 -7622 592650 -7066
rect -8726 -7654 592650 -7622
use user_proj_example  mprj
timestamp 1635497614
transform 1 0 235000 0 1 338000
box 110 0 179846 120000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 4 analog_io[0]
port 1 nsew
rlabel metal2 s 446098 703520 446210 704960 4 analog_io[10]
port 2 nsew
rlabel metal2 s 381146 703520 381258 704960 4 analog_io[11]
port 3 nsew
rlabel metal2 s 316286 703520 316398 704960 4 analog_io[12]
port 4 nsew
rlabel metal2 s 251426 703520 251538 704960 4 analog_io[13]
port 5 nsew
rlabel metal2 s 186474 703520 186586 704960 4 analog_io[14]
port 6 nsew
rlabel metal2 s 121614 703520 121726 704960 4 analog_io[15]
port 7 nsew
rlabel metal2 s 56754 703520 56866 704960 4 analog_io[16]
port 8 nsew
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 9 nsew
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 10 nsew
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 11 nsew
rlabel metal3 s 583520 338452 584960 338692 4 analog_io[1]
port 12 nsew
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 13 nsew
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 14 nsew
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 15 nsew
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 16 nsew
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 17 nsew
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 18 nsew
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 19 nsew
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 20 nsew
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 21 nsew
rlabel metal3 s 583520 391628 584960 391868 4 analog_io[2]
port 22 nsew
rlabel metal3 s 583520 444668 584960 444908 4 analog_io[3]
port 23 nsew
rlabel metal3 s 583520 497844 584960 498084 4 analog_io[4]
port 24 nsew
rlabel metal3 s 583520 551020 584960 551260 4 analog_io[5]
port 25 nsew
rlabel metal3 s 583520 604060 584960 604300 4 analog_io[6]
port 26 nsew
rlabel metal3 s 583520 657236 584960 657476 4 analog_io[7]
port 27 nsew
rlabel metal2 s 575818 703520 575930 704960 4 analog_io[8]
port 28 nsew
rlabel metal2 s 510958 703520 511070 704960 4 analog_io[9]
port 29 nsew
rlabel metal3 s 583520 6476 584960 6716 4 io_in[0]
port 30 nsew
rlabel metal3 s 583520 457996 584960 458236 4 io_in[10]
port 31 nsew
rlabel metal3 s 583520 511172 584960 511412 4 io_in[11]
port 32 nsew
rlabel metal3 s 583520 564212 584960 564452 4 io_in[12]
port 33 nsew
rlabel metal3 s 583520 617388 584960 617628 4 io_in[13]
port 34 nsew
rlabel metal3 s 583520 670564 584960 670804 4 io_in[14]
port 35 nsew
rlabel metal2 s 559626 703520 559738 704960 4 io_in[15]
port 36 nsew
rlabel metal2 s 494766 703520 494878 704960 4 io_in[16]
port 37 nsew
rlabel metal2 s 429814 703520 429926 704960 4 io_in[17]
port 38 nsew
rlabel metal2 s 364954 703520 365066 704960 4 io_in[18]
port 39 nsew
rlabel metal2 s 300094 703520 300206 704960 4 io_in[19]
port 40 nsew
rlabel metal3 s 583520 46188 584960 46428 4 io_in[1]
port 41 nsew
rlabel metal2 s 235142 703520 235254 704960 4 io_in[20]
port 42 nsew
rlabel metal2 s 170282 703520 170394 704960 4 io_in[21]
port 43 nsew
rlabel metal2 s 105422 703520 105534 704960 4 io_in[22]
port 44 nsew
rlabel metal2 s 40470 703520 40582 704960 4 io_in[23]
port 45 nsew
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 46 nsew
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 47 nsew
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 48 nsew
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 49 nsew
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 50 nsew
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 51 nsew
rlabel metal3 s 583520 86036 584960 86276 4 io_in[2]
port 52 nsew
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 53 nsew
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 54 nsew
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 55 nsew
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 56 nsew
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 57 nsew
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 58 nsew
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 59 nsew
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 60 nsew
rlabel metal3 s 583520 125884 584960 126124 4 io_in[3]
port 61 nsew
rlabel metal3 s 583520 165732 584960 165972 4 io_in[4]
port 62 nsew
rlabel metal3 s 583520 205580 584960 205820 4 io_in[5]
port 63 nsew
rlabel metal3 s 583520 245428 584960 245668 4 io_in[6]
port 64 nsew
rlabel metal3 s 583520 298604 584960 298844 4 io_in[7]
port 65 nsew
rlabel metal3 s 583520 351780 584960 352020 4 io_in[8]
port 66 nsew
rlabel metal3 s 583520 404820 584960 405060 4 io_in[9]
port 67 nsew
rlabel metal3 s 583520 32996 584960 33236 4 io_oeb[0]
port 68 nsew
rlabel metal3 s 583520 484516 584960 484756 4 io_oeb[10]
port 69 nsew
rlabel metal3 s 583520 537692 584960 537932 4 io_oeb[11]
port 70 nsew
rlabel metal3 s 583520 590868 584960 591108 4 io_oeb[12]
port 71 nsew
rlabel metal3 s 583520 643908 584960 644148 4 io_oeb[13]
port 72 nsew
rlabel metal3 s 583520 697084 584960 697324 4 io_oeb[14]
port 73 nsew
rlabel metal2 s 527150 703520 527262 704960 4 io_oeb[15]
port 74 nsew
rlabel metal2 s 462290 703520 462402 704960 4 io_oeb[16]
port 75 nsew
rlabel metal2 s 397430 703520 397542 704960 4 io_oeb[17]
port 76 nsew
rlabel metal2 s 332478 703520 332590 704960 4 io_oeb[18]
port 77 nsew
rlabel metal2 s 267618 703520 267730 704960 4 io_oeb[19]
port 78 nsew
rlabel metal3 s 583520 72844 584960 73084 4 io_oeb[1]
port 79 nsew
rlabel metal2 s 202758 703520 202870 704960 4 io_oeb[20]
port 80 nsew
rlabel metal2 s 137806 703520 137918 704960 4 io_oeb[21]
port 81 nsew
rlabel metal2 s 72946 703520 73058 704960 4 io_oeb[22]
port 82 nsew
rlabel metal2 s 8086 703520 8198 704960 4 io_oeb[23]
port 83 nsew
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 84 nsew
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 85 nsew
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 86 nsew
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 87 nsew
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 88 nsew
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 89 nsew
rlabel metal3 s 583520 112692 584960 112932 4 io_oeb[2]
port 90 nsew
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 91 nsew
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 92 nsew
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 93 nsew
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 94 nsew
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 95 nsew
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 96 nsew
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 97 nsew
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 98 nsew
rlabel metal3 s 583520 152540 584960 152780 4 io_oeb[3]
port 99 nsew
rlabel metal3 s 583520 192388 584960 192628 4 io_oeb[4]
port 100 nsew
rlabel metal3 s 583520 232236 584960 232476 4 io_oeb[5]
port 101 nsew
rlabel metal3 s 583520 272084 584960 272324 4 io_oeb[6]
port 102 nsew
rlabel metal3 s 583520 325124 584960 325364 4 io_oeb[7]
port 103 nsew
rlabel metal3 s 583520 378300 584960 378540 4 io_oeb[8]
port 104 nsew
rlabel metal3 s 583520 431476 584960 431716 4 io_oeb[9]
port 105 nsew
rlabel metal3 s 583520 19668 584960 19908 4 io_out[0]
port 106 nsew
rlabel metal3 s 583520 471324 584960 471564 4 io_out[10]
port 107 nsew
rlabel metal3 s 583520 524364 584960 524604 4 io_out[11]
port 108 nsew
rlabel metal3 s 583520 577540 584960 577780 4 io_out[12]
port 109 nsew
rlabel metal3 s 583520 630716 584960 630956 4 io_out[13]
port 110 nsew
rlabel metal3 s 583520 683756 584960 683996 4 io_out[14]
port 111 nsew
rlabel metal2 s 543434 703520 543546 704960 4 io_out[15]
port 112 nsew
rlabel metal2 s 478482 703520 478594 704960 4 io_out[16]
port 113 nsew
rlabel metal2 s 413622 703520 413734 704960 4 io_out[17]
port 114 nsew
rlabel metal2 s 348762 703520 348874 704960 4 io_out[18]
port 115 nsew
rlabel metal2 s 283810 703520 283922 704960 4 io_out[19]
port 116 nsew
rlabel metal3 s 583520 59516 584960 59756 4 io_out[1]
port 117 nsew
rlabel metal2 s 218950 703520 219062 704960 4 io_out[20]
port 118 nsew
rlabel metal2 s 154090 703520 154202 704960 4 io_out[21]
port 119 nsew
rlabel metal2 s 89138 703520 89250 704960 4 io_out[22]
port 120 nsew
rlabel metal2 s 24278 703520 24390 704960 4 io_out[23]
port 121 nsew
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 122 nsew
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 123 nsew
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 124 nsew
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 125 nsew
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 126 nsew
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 127 nsew
rlabel metal3 s 583520 99364 584960 99604 4 io_out[2]
port 128 nsew
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 129 nsew
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 130 nsew
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 131 nsew
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 132 nsew
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 133 nsew
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 134 nsew
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 135 nsew
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 136 nsew
rlabel metal3 s 583520 139212 584960 139452 4 io_out[3]
port 137 nsew
rlabel metal3 s 583520 179060 584960 179300 4 io_out[4]
port 138 nsew
rlabel metal3 s 583520 218908 584960 219148 4 io_out[5]
port 139 nsew
rlabel metal3 s 583520 258756 584960 258996 4 io_out[6]
port 140 nsew
rlabel metal3 s 583520 311932 584960 312172 4 io_out[7]
port 141 nsew
rlabel metal3 s 583520 364972 584960 365212 4 io_out[8]
port 142 nsew
rlabel metal3 s 583520 418148 584960 418388 4 io_out[9]
port 143 nsew
rlabel metal2 s 125846 -960 125958 480 4 la_data_in[0]
port 144 nsew
rlabel metal2 s 480506 -960 480618 480 4 la_data_in[100]
port 145 nsew
rlabel metal2 s 484002 -960 484114 480 4 la_data_in[101]
port 146 nsew
rlabel metal2 s 487590 -960 487702 480 4 la_data_in[102]
port 147 nsew
rlabel metal2 s 491086 -960 491198 480 4 la_data_in[103]
port 148 nsew
rlabel metal2 s 494674 -960 494786 480 4 la_data_in[104]
port 149 nsew
rlabel metal2 s 498170 -960 498282 480 4 la_data_in[105]
port 150 nsew
rlabel metal2 s 501758 -960 501870 480 4 la_data_in[106]
port 151 nsew
rlabel metal2 s 505346 -960 505458 480 4 la_data_in[107]
port 152 nsew
rlabel metal2 s 508842 -960 508954 480 4 la_data_in[108]
port 153 nsew
rlabel metal2 s 512430 -960 512542 480 4 la_data_in[109]
port 154 nsew
rlabel metal2 s 161266 -960 161378 480 4 la_data_in[10]
port 155 nsew
rlabel metal2 s 515926 -960 516038 480 4 la_data_in[110]
port 156 nsew
rlabel metal2 s 519514 -960 519626 480 4 la_data_in[111]
port 157 nsew
rlabel metal2 s 523010 -960 523122 480 4 la_data_in[112]
port 158 nsew
rlabel metal2 s 526598 -960 526710 480 4 la_data_in[113]
port 159 nsew
rlabel metal2 s 530094 -960 530206 480 4 la_data_in[114]
port 160 nsew
rlabel metal2 s 533682 -960 533794 480 4 la_data_in[115]
port 161 nsew
rlabel metal2 s 537178 -960 537290 480 4 la_data_in[116]
port 162 nsew
rlabel metal2 s 540766 -960 540878 480 4 la_data_in[117]
port 163 nsew
rlabel metal2 s 544354 -960 544466 480 4 la_data_in[118]
port 164 nsew
rlabel metal2 s 547850 -960 547962 480 4 la_data_in[119]
port 165 nsew
rlabel metal2 s 164854 -960 164966 480 4 la_data_in[11]
port 166 nsew
rlabel metal2 s 551438 -960 551550 480 4 la_data_in[120]
port 167 nsew
rlabel metal2 s 554934 -960 555046 480 4 la_data_in[121]
port 168 nsew
rlabel metal2 s 558522 -960 558634 480 4 la_data_in[122]
port 169 nsew
rlabel metal2 s 562018 -960 562130 480 4 la_data_in[123]
port 170 nsew
rlabel metal2 s 565606 -960 565718 480 4 la_data_in[124]
port 171 nsew
rlabel metal2 s 569102 -960 569214 480 4 la_data_in[125]
port 172 nsew
rlabel metal2 s 572690 -960 572802 480 4 la_data_in[126]
port 173 nsew
rlabel metal2 s 576278 -960 576390 480 4 la_data_in[127]
port 174 nsew
rlabel metal2 s 168350 -960 168462 480 4 la_data_in[12]
port 175 nsew
rlabel metal2 s 171938 -960 172050 480 4 la_data_in[13]
port 176 nsew
rlabel metal2 s 175434 -960 175546 480 4 la_data_in[14]
port 177 nsew
rlabel metal2 s 179022 -960 179134 480 4 la_data_in[15]
port 178 nsew
rlabel metal2 s 182518 -960 182630 480 4 la_data_in[16]
port 179 nsew
rlabel metal2 s 186106 -960 186218 480 4 la_data_in[17]
port 180 nsew
rlabel metal2 s 189694 -960 189806 480 4 la_data_in[18]
port 181 nsew
rlabel metal2 s 193190 -960 193302 480 4 la_data_in[19]
port 182 nsew
rlabel metal2 s 129342 -960 129454 480 4 la_data_in[1]
port 183 nsew
rlabel metal2 s 196778 -960 196890 480 4 la_data_in[20]
port 184 nsew
rlabel metal2 s 200274 -960 200386 480 4 la_data_in[21]
port 185 nsew
rlabel metal2 s 203862 -960 203974 480 4 la_data_in[22]
port 186 nsew
rlabel metal2 s 207358 -960 207470 480 4 la_data_in[23]
port 187 nsew
rlabel metal2 s 210946 -960 211058 480 4 la_data_in[24]
port 188 nsew
rlabel metal2 s 214442 -960 214554 480 4 la_data_in[25]
port 189 nsew
rlabel metal2 s 218030 -960 218142 480 4 la_data_in[26]
port 190 nsew
rlabel metal2 s 221526 -960 221638 480 4 la_data_in[27]
port 191 nsew
rlabel metal2 s 225114 -960 225226 480 4 la_data_in[28]
port 192 nsew
rlabel metal2 s 228702 -960 228814 480 4 la_data_in[29]
port 193 nsew
rlabel metal2 s 132930 -960 133042 480 4 la_data_in[2]
port 194 nsew
rlabel metal2 s 232198 -960 232310 480 4 la_data_in[30]
port 195 nsew
rlabel metal2 s 235786 -960 235898 480 4 la_data_in[31]
port 196 nsew
rlabel metal2 s 239282 -960 239394 480 4 la_data_in[32]
port 197 nsew
rlabel metal2 s 242870 -960 242982 480 4 la_data_in[33]
port 198 nsew
rlabel metal2 s 246366 -960 246478 480 4 la_data_in[34]
port 199 nsew
rlabel metal2 s 249954 -960 250066 480 4 la_data_in[35]
port 200 nsew
rlabel metal2 s 253450 -960 253562 480 4 la_data_in[36]
port 201 nsew
rlabel metal2 s 257038 -960 257150 480 4 la_data_in[37]
port 202 nsew
rlabel metal2 s 260626 -960 260738 480 4 la_data_in[38]
port 203 nsew
rlabel metal2 s 264122 -960 264234 480 4 la_data_in[39]
port 204 nsew
rlabel metal2 s 136426 -960 136538 480 4 la_data_in[3]
port 205 nsew
rlabel metal2 s 267710 -960 267822 480 4 la_data_in[40]
port 206 nsew
rlabel metal2 s 271206 -960 271318 480 4 la_data_in[41]
port 207 nsew
rlabel metal2 s 274794 -960 274906 480 4 la_data_in[42]
port 208 nsew
rlabel metal2 s 278290 -960 278402 480 4 la_data_in[43]
port 209 nsew
rlabel metal2 s 281878 -960 281990 480 4 la_data_in[44]
port 210 nsew
rlabel metal2 s 285374 -960 285486 480 4 la_data_in[45]
port 211 nsew
rlabel metal2 s 288962 -960 289074 480 4 la_data_in[46]
port 212 nsew
rlabel metal2 s 292550 -960 292662 480 4 la_data_in[47]
port 213 nsew
rlabel metal2 s 296046 -960 296158 480 4 la_data_in[48]
port 214 nsew
rlabel metal2 s 299634 -960 299746 480 4 la_data_in[49]
port 215 nsew
rlabel metal2 s 140014 -960 140126 480 4 la_data_in[4]
port 216 nsew
rlabel metal2 s 303130 -960 303242 480 4 la_data_in[50]
port 217 nsew
rlabel metal2 s 306718 -960 306830 480 4 la_data_in[51]
port 218 nsew
rlabel metal2 s 310214 -960 310326 480 4 la_data_in[52]
port 219 nsew
rlabel metal2 s 313802 -960 313914 480 4 la_data_in[53]
port 220 nsew
rlabel metal2 s 317298 -960 317410 480 4 la_data_in[54]
port 221 nsew
rlabel metal2 s 320886 -960 320998 480 4 la_data_in[55]
port 222 nsew
rlabel metal2 s 324382 -960 324494 480 4 la_data_in[56]
port 223 nsew
rlabel metal2 s 327970 -960 328082 480 4 la_data_in[57]
port 224 nsew
rlabel metal2 s 331558 -960 331670 480 4 la_data_in[58]
port 225 nsew
rlabel metal2 s 335054 -960 335166 480 4 la_data_in[59]
port 226 nsew
rlabel metal2 s 143510 -960 143622 480 4 la_data_in[5]
port 227 nsew
rlabel metal2 s 338642 -960 338754 480 4 la_data_in[60]
port 228 nsew
rlabel metal2 s 342138 -960 342250 480 4 la_data_in[61]
port 229 nsew
rlabel metal2 s 345726 -960 345838 480 4 la_data_in[62]
port 230 nsew
rlabel metal2 s 349222 -960 349334 480 4 la_data_in[63]
port 231 nsew
rlabel metal2 s 352810 -960 352922 480 4 la_data_in[64]
port 232 nsew
rlabel metal2 s 356306 -960 356418 480 4 la_data_in[65]
port 233 nsew
rlabel metal2 s 359894 -960 360006 480 4 la_data_in[66]
port 234 nsew
rlabel metal2 s 363482 -960 363594 480 4 la_data_in[67]
port 235 nsew
rlabel metal2 s 366978 -960 367090 480 4 la_data_in[68]
port 236 nsew
rlabel metal2 s 370566 -960 370678 480 4 la_data_in[69]
port 237 nsew
rlabel metal2 s 147098 -960 147210 480 4 la_data_in[6]
port 238 nsew
rlabel metal2 s 374062 -960 374174 480 4 la_data_in[70]
port 239 nsew
rlabel metal2 s 377650 -960 377762 480 4 la_data_in[71]
port 240 nsew
rlabel metal2 s 381146 -960 381258 480 4 la_data_in[72]
port 241 nsew
rlabel metal2 s 384734 -960 384846 480 4 la_data_in[73]
port 242 nsew
rlabel metal2 s 388230 -960 388342 480 4 la_data_in[74]
port 243 nsew
rlabel metal2 s 391818 -960 391930 480 4 la_data_in[75]
port 244 nsew
rlabel metal2 s 395314 -960 395426 480 4 la_data_in[76]
port 245 nsew
rlabel metal2 s 398902 -960 399014 480 4 la_data_in[77]
port 246 nsew
rlabel metal2 s 402490 -960 402602 480 4 la_data_in[78]
port 247 nsew
rlabel metal2 s 405986 -960 406098 480 4 la_data_in[79]
port 248 nsew
rlabel metal2 s 150594 -960 150706 480 4 la_data_in[7]
port 249 nsew
rlabel metal2 s 409574 -960 409686 480 4 la_data_in[80]
port 250 nsew
rlabel metal2 s 413070 -960 413182 480 4 la_data_in[81]
port 251 nsew
rlabel metal2 s 416658 -960 416770 480 4 la_data_in[82]
port 252 nsew
rlabel metal2 s 420154 -960 420266 480 4 la_data_in[83]
port 253 nsew
rlabel metal2 s 423742 -960 423854 480 4 la_data_in[84]
port 254 nsew
rlabel metal2 s 427238 -960 427350 480 4 la_data_in[85]
port 255 nsew
rlabel metal2 s 430826 -960 430938 480 4 la_data_in[86]
port 256 nsew
rlabel metal2 s 434414 -960 434526 480 4 la_data_in[87]
port 257 nsew
rlabel metal2 s 437910 -960 438022 480 4 la_data_in[88]
port 258 nsew
rlabel metal2 s 441498 -960 441610 480 4 la_data_in[89]
port 259 nsew
rlabel metal2 s 154182 -960 154294 480 4 la_data_in[8]
port 260 nsew
rlabel metal2 s 444994 -960 445106 480 4 la_data_in[90]
port 261 nsew
rlabel metal2 s 448582 -960 448694 480 4 la_data_in[91]
port 262 nsew
rlabel metal2 s 452078 -960 452190 480 4 la_data_in[92]
port 263 nsew
rlabel metal2 s 455666 -960 455778 480 4 la_data_in[93]
port 264 nsew
rlabel metal2 s 459162 -960 459274 480 4 la_data_in[94]
port 265 nsew
rlabel metal2 s 462750 -960 462862 480 4 la_data_in[95]
port 266 nsew
rlabel metal2 s 466246 -960 466358 480 4 la_data_in[96]
port 267 nsew
rlabel metal2 s 469834 -960 469946 480 4 la_data_in[97]
port 268 nsew
rlabel metal2 s 473422 -960 473534 480 4 la_data_in[98]
port 269 nsew
rlabel metal2 s 476918 -960 477030 480 4 la_data_in[99]
port 270 nsew
rlabel metal2 s 157770 -960 157882 480 4 la_data_in[9]
port 271 nsew
rlabel metal2 s 126950 -960 127062 480 4 la_data_out[0]
port 272 nsew
rlabel metal2 s 481702 -960 481814 480 4 la_data_out[100]
port 273 nsew
rlabel metal2 s 485198 -960 485310 480 4 la_data_out[101]
port 274 nsew
rlabel metal2 s 488786 -960 488898 480 4 la_data_out[102]
port 275 nsew
rlabel metal2 s 492282 -960 492394 480 4 la_data_out[103]
port 276 nsew
rlabel metal2 s 495870 -960 495982 480 4 la_data_out[104]
port 277 nsew
rlabel metal2 s 499366 -960 499478 480 4 la_data_out[105]
port 278 nsew
rlabel metal2 s 502954 -960 503066 480 4 la_data_out[106]
port 279 nsew
rlabel metal2 s 506450 -960 506562 480 4 la_data_out[107]
port 280 nsew
rlabel metal2 s 510038 -960 510150 480 4 la_data_out[108]
port 281 nsew
rlabel metal2 s 513534 -960 513646 480 4 la_data_out[109]
port 282 nsew
rlabel metal2 s 162462 -960 162574 480 4 la_data_out[10]
port 283 nsew
rlabel metal2 s 517122 -960 517234 480 4 la_data_out[110]
port 284 nsew
rlabel metal2 s 520710 -960 520822 480 4 la_data_out[111]
port 285 nsew
rlabel metal2 s 524206 -960 524318 480 4 la_data_out[112]
port 286 nsew
rlabel metal2 s 527794 -960 527906 480 4 la_data_out[113]
port 287 nsew
rlabel metal2 s 531290 -960 531402 480 4 la_data_out[114]
port 288 nsew
rlabel metal2 s 534878 -960 534990 480 4 la_data_out[115]
port 289 nsew
rlabel metal2 s 538374 -960 538486 480 4 la_data_out[116]
port 290 nsew
rlabel metal2 s 541962 -960 542074 480 4 la_data_out[117]
port 291 nsew
rlabel metal2 s 545458 -960 545570 480 4 la_data_out[118]
port 292 nsew
rlabel metal2 s 549046 -960 549158 480 4 la_data_out[119]
port 293 nsew
rlabel metal2 s 166050 -960 166162 480 4 la_data_out[11]
port 294 nsew
rlabel metal2 s 552634 -960 552746 480 4 la_data_out[120]
port 295 nsew
rlabel metal2 s 556130 -960 556242 480 4 la_data_out[121]
port 296 nsew
rlabel metal2 s 559718 -960 559830 480 4 la_data_out[122]
port 297 nsew
rlabel metal2 s 563214 -960 563326 480 4 la_data_out[123]
port 298 nsew
rlabel metal2 s 566802 -960 566914 480 4 la_data_out[124]
port 299 nsew
rlabel metal2 s 570298 -960 570410 480 4 la_data_out[125]
port 300 nsew
rlabel metal2 s 573886 -960 573998 480 4 la_data_out[126]
port 301 nsew
rlabel metal2 s 577382 -960 577494 480 4 la_data_out[127]
port 302 nsew
rlabel metal2 s 169546 -960 169658 480 4 la_data_out[12]
port 303 nsew
rlabel metal2 s 173134 -960 173246 480 4 la_data_out[13]
port 304 nsew
rlabel metal2 s 176630 -960 176742 480 4 la_data_out[14]
port 305 nsew
rlabel metal2 s 180218 -960 180330 480 4 la_data_out[15]
port 306 nsew
rlabel metal2 s 183714 -960 183826 480 4 la_data_out[16]
port 307 nsew
rlabel metal2 s 187302 -960 187414 480 4 la_data_out[17]
port 308 nsew
rlabel metal2 s 190798 -960 190910 480 4 la_data_out[18]
port 309 nsew
rlabel metal2 s 194386 -960 194498 480 4 la_data_out[19]
port 310 nsew
rlabel metal2 s 130538 -960 130650 480 4 la_data_out[1]
port 311 nsew
rlabel metal2 s 197882 -960 197994 480 4 la_data_out[20]
port 312 nsew
rlabel metal2 s 201470 -960 201582 480 4 la_data_out[21]
port 313 nsew
rlabel metal2 s 205058 -960 205170 480 4 la_data_out[22]
port 314 nsew
rlabel metal2 s 208554 -960 208666 480 4 la_data_out[23]
port 315 nsew
rlabel metal2 s 212142 -960 212254 480 4 la_data_out[24]
port 316 nsew
rlabel metal2 s 215638 -960 215750 480 4 la_data_out[25]
port 317 nsew
rlabel metal2 s 219226 -960 219338 480 4 la_data_out[26]
port 318 nsew
rlabel metal2 s 222722 -960 222834 480 4 la_data_out[27]
port 319 nsew
rlabel metal2 s 226310 -960 226422 480 4 la_data_out[28]
port 320 nsew
rlabel metal2 s 229806 -960 229918 480 4 la_data_out[29]
port 321 nsew
rlabel metal2 s 134126 -960 134238 480 4 la_data_out[2]
port 322 nsew
rlabel metal2 s 233394 -960 233506 480 4 la_data_out[30]
port 323 nsew
rlabel metal2 s 236982 -960 237094 480 4 la_data_out[31]
port 324 nsew
rlabel metal2 s 240478 -960 240590 480 4 la_data_out[32]
port 325 nsew
rlabel metal2 s 244066 -960 244178 480 4 la_data_out[33]
port 326 nsew
rlabel metal2 s 247562 -960 247674 480 4 la_data_out[34]
port 327 nsew
rlabel metal2 s 251150 -960 251262 480 4 la_data_out[35]
port 328 nsew
rlabel metal2 s 254646 -960 254758 480 4 la_data_out[36]
port 329 nsew
rlabel metal2 s 258234 -960 258346 480 4 la_data_out[37]
port 330 nsew
rlabel metal2 s 261730 -960 261842 480 4 la_data_out[38]
port 331 nsew
rlabel metal2 s 265318 -960 265430 480 4 la_data_out[39]
port 332 nsew
rlabel metal2 s 137622 -960 137734 480 4 la_data_out[3]
port 333 nsew
rlabel metal2 s 268814 -960 268926 480 4 la_data_out[40]
port 334 nsew
rlabel metal2 s 272402 -960 272514 480 4 la_data_out[41]
port 335 nsew
rlabel metal2 s 275990 -960 276102 480 4 la_data_out[42]
port 336 nsew
rlabel metal2 s 279486 -960 279598 480 4 la_data_out[43]
port 337 nsew
rlabel metal2 s 283074 -960 283186 480 4 la_data_out[44]
port 338 nsew
rlabel metal2 s 286570 -960 286682 480 4 la_data_out[45]
port 339 nsew
rlabel metal2 s 290158 -960 290270 480 4 la_data_out[46]
port 340 nsew
rlabel metal2 s 293654 -960 293766 480 4 la_data_out[47]
port 341 nsew
rlabel metal2 s 297242 -960 297354 480 4 la_data_out[48]
port 342 nsew
rlabel metal2 s 300738 -960 300850 480 4 la_data_out[49]
port 343 nsew
rlabel metal2 s 141210 -960 141322 480 4 la_data_out[4]
port 344 nsew
rlabel metal2 s 304326 -960 304438 480 4 la_data_out[50]
port 345 nsew
rlabel metal2 s 307914 -960 308026 480 4 la_data_out[51]
port 346 nsew
rlabel metal2 s 311410 -960 311522 480 4 la_data_out[52]
port 347 nsew
rlabel metal2 s 314998 -960 315110 480 4 la_data_out[53]
port 348 nsew
rlabel metal2 s 318494 -960 318606 480 4 la_data_out[54]
port 349 nsew
rlabel metal2 s 322082 -960 322194 480 4 la_data_out[55]
port 350 nsew
rlabel metal2 s 325578 -960 325690 480 4 la_data_out[56]
port 351 nsew
rlabel metal2 s 329166 -960 329278 480 4 la_data_out[57]
port 352 nsew
rlabel metal2 s 332662 -960 332774 480 4 la_data_out[58]
port 353 nsew
rlabel metal2 s 336250 -960 336362 480 4 la_data_out[59]
port 354 nsew
rlabel metal2 s 144706 -960 144818 480 4 la_data_out[5]
port 355 nsew
rlabel metal2 s 339838 -960 339950 480 4 la_data_out[60]
port 356 nsew
rlabel metal2 s 343334 -960 343446 480 4 la_data_out[61]
port 357 nsew
rlabel metal2 s 346922 -960 347034 480 4 la_data_out[62]
port 358 nsew
rlabel metal2 s 350418 -960 350530 480 4 la_data_out[63]
port 359 nsew
rlabel metal2 s 354006 -960 354118 480 4 la_data_out[64]
port 360 nsew
rlabel metal2 s 357502 -960 357614 480 4 la_data_out[65]
port 361 nsew
rlabel metal2 s 361090 -960 361202 480 4 la_data_out[66]
port 362 nsew
rlabel metal2 s 364586 -960 364698 480 4 la_data_out[67]
port 363 nsew
rlabel metal2 s 368174 -960 368286 480 4 la_data_out[68]
port 364 nsew
rlabel metal2 s 371670 -960 371782 480 4 la_data_out[69]
port 365 nsew
rlabel metal2 s 148294 -960 148406 480 4 la_data_out[6]
port 366 nsew
rlabel metal2 s 375258 -960 375370 480 4 la_data_out[70]
port 367 nsew
rlabel metal2 s 378846 -960 378958 480 4 la_data_out[71]
port 368 nsew
rlabel metal2 s 382342 -960 382454 480 4 la_data_out[72]
port 369 nsew
rlabel metal2 s 385930 -960 386042 480 4 la_data_out[73]
port 370 nsew
rlabel metal2 s 389426 -960 389538 480 4 la_data_out[74]
port 371 nsew
rlabel metal2 s 393014 -960 393126 480 4 la_data_out[75]
port 372 nsew
rlabel metal2 s 396510 -960 396622 480 4 la_data_out[76]
port 373 nsew
rlabel metal2 s 400098 -960 400210 480 4 la_data_out[77]
port 374 nsew
rlabel metal2 s 403594 -960 403706 480 4 la_data_out[78]
port 375 nsew
rlabel metal2 s 407182 -960 407294 480 4 la_data_out[79]
port 376 nsew
rlabel metal2 s 151790 -960 151902 480 4 la_data_out[7]
port 377 nsew
rlabel metal2 s 410770 -960 410882 480 4 la_data_out[80]
port 378 nsew
rlabel metal2 s 414266 -960 414378 480 4 la_data_out[81]
port 379 nsew
rlabel metal2 s 417854 -960 417966 480 4 la_data_out[82]
port 380 nsew
rlabel metal2 s 421350 -960 421462 480 4 la_data_out[83]
port 381 nsew
rlabel metal2 s 424938 -960 425050 480 4 la_data_out[84]
port 382 nsew
rlabel metal2 s 428434 -960 428546 480 4 la_data_out[85]
port 383 nsew
rlabel metal2 s 432022 -960 432134 480 4 la_data_out[86]
port 384 nsew
rlabel metal2 s 435518 -960 435630 480 4 la_data_out[87]
port 385 nsew
rlabel metal2 s 439106 -960 439218 480 4 la_data_out[88]
port 386 nsew
rlabel metal2 s 442602 -960 442714 480 4 la_data_out[89]
port 387 nsew
rlabel metal2 s 155378 -960 155490 480 4 la_data_out[8]
port 388 nsew
rlabel metal2 s 446190 -960 446302 480 4 la_data_out[90]
port 389 nsew
rlabel metal2 s 449778 -960 449890 480 4 la_data_out[91]
port 390 nsew
rlabel metal2 s 453274 -960 453386 480 4 la_data_out[92]
port 391 nsew
rlabel metal2 s 456862 -960 456974 480 4 la_data_out[93]
port 392 nsew
rlabel metal2 s 460358 -960 460470 480 4 la_data_out[94]
port 393 nsew
rlabel metal2 s 463946 -960 464058 480 4 la_data_out[95]
port 394 nsew
rlabel metal2 s 467442 -960 467554 480 4 la_data_out[96]
port 395 nsew
rlabel metal2 s 471030 -960 471142 480 4 la_data_out[97]
port 396 nsew
rlabel metal2 s 474526 -960 474638 480 4 la_data_out[98]
port 397 nsew
rlabel metal2 s 478114 -960 478226 480 4 la_data_out[99]
port 398 nsew
rlabel metal2 s 158874 -960 158986 480 4 la_data_out[9]
port 399 nsew
rlabel metal2 s 128146 -960 128258 480 4 la_oenb[0]
port 400 nsew
rlabel metal2 s 482806 -960 482918 480 4 la_oenb[100]
port 401 nsew
rlabel metal2 s 486394 -960 486506 480 4 la_oenb[101]
port 402 nsew
rlabel metal2 s 489890 -960 490002 480 4 la_oenb[102]
port 403 nsew
rlabel metal2 s 493478 -960 493590 480 4 la_oenb[103]
port 404 nsew
rlabel metal2 s 497066 -960 497178 480 4 la_oenb[104]
port 405 nsew
rlabel metal2 s 500562 -960 500674 480 4 la_oenb[105]
port 406 nsew
rlabel metal2 s 504150 -960 504262 480 4 la_oenb[106]
port 407 nsew
rlabel metal2 s 507646 -960 507758 480 4 la_oenb[107]
port 408 nsew
rlabel metal2 s 511234 -960 511346 480 4 la_oenb[108]
port 409 nsew
rlabel metal2 s 514730 -960 514842 480 4 la_oenb[109]
port 410 nsew
rlabel metal2 s 163658 -960 163770 480 4 la_oenb[10]
port 411 nsew
rlabel metal2 s 518318 -960 518430 480 4 la_oenb[110]
port 412 nsew
rlabel metal2 s 521814 -960 521926 480 4 la_oenb[111]
port 413 nsew
rlabel metal2 s 525402 -960 525514 480 4 la_oenb[112]
port 414 nsew
rlabel metal2 s 528990 -960 529102 480 4 la_oenb[113]
port 415 nsew
rlabel metal2 s 532486 -960 532598 480 4 la_oenb[114]
port 416 nsew
rlabel metal2 s 536074 -960 536186 480 4 la_oenb[115]
port 417 nsew
rlabel metal2 s 539570 -960 539682 480 4 la_oenb[116]
port 418 nsew
rlabel metal2 s 543158 -960 543270 480 4 la_oenb[117]
port 419 nsew
rlabel metal2 s 546654 -960 546766 480 4 la_oenb[118]
port 420 nsew
rlabel metal2 s 550242 -960 550354 480 4 la_oenb[119]
port 421 nsew
rlabel metal2 s 167154 -960 167266 480 4 la_oenb[11]
port 422 nsew
rlabel metal2 s 553738 -960 553850 480 4 la_oenb[120]
port 423 nsew
rlabel metal2 s 557326 -960 557438 480 4 la_oenb[121]
port 424 nsew
rlabel metal2 s 560822 -960 560934 480 4 la_oenb[122]
port 425 nsew
rlabel metal2 s 564410 -960 564522 480 4 la_oenb[123]
port 426 nsew
rlabel metal2 s 567998 -960 568110 480 4 la_oenb[124]
port 427 nsew
rlabel metal2 s 571494 -960 571606 480 4 la_oenb[125]
port 428 nsew
rlabel metal2 s 575082 -960 575194 480 4 la_oenb[126]
port 429 nsew
rlabel metal2 s 578578 -960 578690 480 4 la_oenb[127]
port 430 nsew
rlabel metal2 s 170742 -960 170854 480 4 la_oenb[12]
port 431 nsew
rlabel metal2 s 174238 -960 174350 480 4 la_oenb[13]
port 432 nsew
rlabel metal2 s 177826 -960 177938 480 4 la_oenb[14]
port 433 nsew
rlabel metal2 s 181414 -960 181526 480 4 la_oenb[15]
port 434 nsew
rlabel metal2 s 184910 -960 185022 480 4 la_oenb[16]
port 435 nsew
rlabel metal2 s 188498 -960 188610 480 4 la_oenb[17]
port 436 nsew
rlabel metal2 s 191994 -960 192106 480 4 la_oenb[18]
port 437 nsew
rlabel metal2 s 195582 -960 195694 480 4 la_oenb[19]
port 438 nsew
rlabel metal2 s 131734 -960 131846 480 4 la_oenb[1]
port 439 nsew
rlabel metal2 s 199078 -960 199190 480 4 la_oenb[20]
port 440 nsew
rlabel metal2 s 202666 -960 202778 480 4 la_oenb[21]
port 441 nsew
rlabel metal2 s 206162 -960 206274 480 4 la_oenb[22]
port 442 nsew
rlabel metal2 s 209750 -960 209862 480 4 la_oenb[23]
port 443 nsew
rlabel metal2 s 213338 -960 213450 480 4 la_oenb[24]
port 444 nsew
rlabel metal2 s 216834 -960 216946 480 4 la_oenb[25]
port 445 nsew
rlabel metal2 s 220422 -960 220534 480 4 la_oenb[26]
port 446 nsew
rlabel metal2 s 223918 -960 224030 480 4 la_oenb[27]
port 447 nsew
rlabel metal2 s 227506 -960 227618 480 4 la_oenb[28]
port 448 nsew
rlabel metal2 s 231002 -960 231114 480 4 la_oenb[29]
port 449 nsew
rlabel metal2 s 135230 -960 135342 480 4 la_oenb[2]
port 450 nsew
rlabel metal2 s 234590 -960 234702 480 4 la_oenb[30]
port 451 nsew
rlabel metal2 s 238086 -960 238198 480 4 la_oenb[31]
port 452 nsew
rlabel metal2 s 241674 -960 241786 480 4 la_oenb[32]
port 453 nsew
rlabel metal2 s 245170 -960 245282 480 4 la_oenb[33]
port 454 nsew
rlabel metal2 s 248758 -960 248870 480 4 la_oenb[34]
port 455 nsew
rlabel metal2 s 252346 -960 252458 480 4 la_oenb[35]
port 456 nsew
rlabel metal2 s 255842 -960 255954 480 4 la_oenb[36]
port 457 nsew
rlabel metal2 s 259430 -960 259542 480 4 la_oenb[37]
port 458 nsew
rlabel metal2 s 262926 -960 263038 480 4 la_oenb[38]
port 459 nsew
rlabel metal2 s 266514 -960 266626 480 4 la_oenb[39]
port 460 nsew
rlabel metal2 s 138818 -960 138930 480 4 la_oenb[3]
port 461 nsew
rlabel metal2 s 270010 -960 270122 480 4 la_oenb[40]
port 462 nsew
rlabel metal2 s 273598 -960 273710 480 4 la_oenb[41]
port 463 nsew
rlabel metal2 s 277094 -960 277206 480 4 la_oenb[42]
port 464 nsew
rlabel metal2 s 280682 -960 280794 480 4 la_oenb[43]
port 465 nsew
rlabel metal2 s 284270 -960 284382 480 4 la_oenb[44]
port 466 nsew
rlabel metal2 s 287766 -960 287878 480 4 la_oenb[45]
port 467 nsew
rlabel metal2 s 291354 -960 291466 480 4 la_oenb[46]
port 468 nsew
rlabel metal2 s 294850 -960 294962 480 4 la_oenb[47]
port 469 nsew
rlabel metal2 s 298438 -960 298550 480 4 la_oenb[48]
port 470 nsew
rlabel metal2 s 301934 -960 302046 480 4 la_oenb[49]
port 471 nsew
rlabel metal2 s 142406 -960 142518 480 4 la_oenb[4]
port 472 nsew
rlabel metal2 s 305522 -960 305634 480 4 la_oenb[50]
port 473 nsew
rlabel metal2 s 309018 -960 309130 480 4 la_oenb[51]
port 474 nsew
rlabel metal2 s 312606 -960 312718 480 4 la_oenb[52]
port 475 nsew
rlabel metal2 s 316194 -960 316306 480 4 la_oenb[53]
port 476 nsew
rlabel metal2 s 319690 -960 319802 480 4 la_oenb[54]
port 477 nsew
rlabel metal2 s 323278 -960 323390 480 4 la_oenb[55]
port 478 nsew
rlabel metal2 s 326774 -960 326886 480 4 la_oenb[56]
port 479 nsew
rlabel metal2 s 330362 -960 330474 480 4 la_oenb[57]
port 480 nsew
rlabel metal2 s 333858 -960 333970 480 4 la_oenb[58]
port 481 nsew
rlabel metal2 s 337446 -960 337558 480 4 la_oenb[59]
port 482 nsew
rlabel metal2 s 145902 -960 146014 480 4 la_oenb[5]
port 483 nsew
rlabel metal2 s 340942 -960 341054 480 4 la_oenb[60]
port 484 nsew
rlabel metal2 s 344530 -960 344642 480 4 la_oenb[61]
port 485 nsew
rlabel metal2 s 348026 -960 348138 480 4 la_oenb[62]
port 486 nsew
rlabel metal2 s 351614 -960 351726 480 4 la_oenb[63]
port 487 nsew
rlabel metal2 s 355202 -960 355314 480 4 la_oenb[64]
port 488 nsew
rlabel metal2 s 358698 -960 358810 480 4 la_oenb[65]
port 489 nsew
rlabel metal2 s 362286 -960 362398 480 4 la_oenb[66]
port 490 nsew
rlabel metal2 s 365782 -960 365894 480 4 la_oenb[67]
port 491 nsew
rlabel metal2 s 369370 -960 369482 480 4 la_oenb[68]
port 492 nsew
rlabel metal2 s 372866 -960 372978 480 4 la_oenb[69]
port 493 nsew
rlabel metal2 s 149490 -960 149602 480 4 la_oenb[6]
port 494 nsew
rlabel metal2 s 376454 -960 376566 480 4 la_oenb[70]
port 495 nsew
rlabel metal2 s 379950 -960 380062 480 4 la_oenb[71]
port 496 nsew
rlabel metal2 s 383538 -960 383650 480 4 la_oenb[72]
port 497 nsew
rlabel metal2 s 387126 -960 387238 480 4 la_oenb[73]
port 498 nsew
rlabel metal2 s 390622 -960 390734 480 4 la_oenb[74]
port 499 nsew
rlabel metal2 s 394210 -960 394322 480 4 la_oenb[75]
port 500 nsew
rlabel metal2 s 397706 -960 397818 480 4 la_oenb[76]
port 501 nsew
rlabel metal2 s 401294 -960 401406 480 4 la_oenb[77]
port 502 nsew
rlabel metal2 s 404790 -960 404902 480 4 la_oenb[78]
port 503 nsew
rlabel metal2 s 408378 -960 408490 480 4 la_oenb[79]
port 504 nsew
rlabel metal2 s 152986 -960 153098 480 4 la_oenb[7]
port 505 nsew
rlabel metal2 s 411874 -960 411986 480 4 la_oenb[80]
port 506 nsew
rlabel metal2 s 415462 -960 415574 480 4 la_oenb[81]
port 507 nsew
rlabel metal2 s 418958 -960 419070 480 4 la_oenb[82]
port 508 nsew
rlabel metal2 s 422546 -960 422658 480 4 la_oenb[83]
port 509 nsew
rlabel metal2 s 426134 -960 426246 480 4 la_oenb[84]
port 510 nsew
rlabel metal2 s 429630 -960 429742 480 4 la_oenb[85]
port 511 nsew
rlabel metal2 s 433218 -960 433330 480 4 la_oenb[86]
port 512 nsew
rlabel metal2 s 436714 -960 436826 480 4 la_oenb[87]
port 513 nsew
rlabel metal2 s 440302 -960 440414 480 4 la_oenb[88]
port 514 nsew
rlabel metal2 s 443798 -960 443910 480 4 la_oenb[89]
port 515 nsew
rlabel metal2 s 156574 -960 156686 480 4 la_oenb[8]
port 516 nsew
rlabel metal2 s 447386 -960 447498 480 4 la_oenb[90]
port 517 nsew
rlabel metal2 s 450882 -960 450994 480 4 la_oenb[91]
port 518 nsew
rlabel metal2 s 454470 -960 454582 480 4 la_oenb[92]
port 519 nsew
rlabel metal2 s 458058 -960 458170 480 4 la_oenb[93]
port 520 nsew
rlabel metal2 s 461554 -960 461666 480 4 la_oenb[94]
port 521 nsew
rlabel metal2 s 465142 -960 465254 480 4 la_oenb[95]
port 522 nsew
rlabel metal2 s 468638 -960 468750 480 4 la_oenb[96]
port 523 nsew
rlabel metal2 s 472226 -960 472338 480 4 la_oenb[97]
port 524 nsew
rlabel metal2 s 475722 -960 475834 480 4 la_oenb[98]
port 525 nsew
rlabel metal2 s 479310 -960 479422 480 4 la_oenb[99]
port 526 nsew
rlabel metal2 s 160070 -960 160182 480 4 la_oenb[9]
port 527 nsew
rlabel metal2 s 579774 -960 579886 480 4 user_clock2
port 528 nsew
rlabel metal2 s 580970 -960 581082 480 4 user_irq[0]
port 529 nsew
rlabel metal2 s 582166 -960 582278 480 4 user_irq[1]
port 530 nsew
rlabel metal2 s 583362 -960 583474 480 4 user_irq[2]
port 531 nsew
rlabel metal5 s -2006 -934 585930 -314 4 vccd1
port 532 nsew
rlabel metal5 s -2966 2866 586890 3486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 38866 586890 39486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 74866 586890 75486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 110866 586890 111486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 146866 586890 147486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 182866 586890 183486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 218866 586890 219486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 254866 586890 255486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 290866 586890 291486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 326866 586890 327486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 362866 586890 363486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 398866 586890 399486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 434866 586890 435486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 470866 586890 471486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 506866 586890 507486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 542866 586890 543486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 578866 586890 579486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 614866 586890 615486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 650866 586890 651486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 686866 586890 687486 4 vccd1
port 532 nsew
rlabel metal5 s -2006 704250 585930 704870 4 vccd1
port 532 nsew
rlabel metal4 s 253794 -1894 254414 338000 4 vccd1
port 532 nsew
rlabel metal4 s 289794 -1894 290414 338000 4 vccd1
port 532 nsew
rlabel metal4 s 325794 -1894 326414 338000 4 vccd1
port 532 nsew
rlabel metal4 s 361794 -1894 362414 338000 4 vccd1
port 532 nsew
rlabel metal4 s 397794 -1894 398414 338000 4 vccd1
port 532 nsew
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 532 nsew
rlabel metal4 s 585310 -934 585930 704870 4 vccd1
port 532 nsew
rlabel metal4 s 1794 -1894 2414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 37794 -1894 38414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 73794 -1894 74414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 109794 -1894 110414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 145794 -1894 146414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 181794 -1894 182414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 217794 -1894 218414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 253794 458000 254414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 289794 458000 290414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 325794 458000 326414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 361794 458000 362414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 397794 458000 398414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 433794 -1894 434414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 469794 -1894 470414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 505794 -1894 506414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 541794 -1894 542414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 577794 -1894 578414 705830 4 vccd1
port 532 nsew
rlabel metal5 s -3926 -2854 587850 -2234 4 vccd2
port 533 nsew
rlabel metal5 s -4886 6586 588810 7206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 42586 588810 43206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 78586 588810 79206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 114586 588810 115206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 150586 588810 151206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 186586 588810 187206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 222586 588810 223206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 258586 588810 259206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 294586 588810 295206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 330586 588810 331206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 366586 588810 367206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 402586 588810 403206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 438586 588810 439206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 474586 588810 475206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 510586 588810 511206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 546586 588810 547206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 582586 588810 583206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 618586 588810 619206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 654586 588810 655206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 690586 588810 691206 4 vccd2
port 533 nsew
rlabel metal5 s -3926 706170 587850 706790 4 vccd2
port 533 nsew
rlabel metal4 s 257514 -3814 258134 336000 4 vccd2
port 533 nsew
rlabel metal4 s 293514 -3814 294134 336000 4 vccd2
port 533 nsew
rlabel metal4 s 329514 -3814 330134 336000 4 vccd2
port 533 nsew
rlabel metal4 s 365514 -3814 366134 336000 4 vccd2
port 533 nsew
rlabel metal4 s 401514 -3814 402134 336000 4 vccd2
port 533 nsew
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 533 nsew
rlabel metal4 s 587230 -2854 587850 706790 4 vccd2
port 533 nsew
rlabel metal4 s 5514 -3814 6134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 41514 -3814 42134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 77514 -3814 78134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 113514 -3814 114134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 149514 -3814 150134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 185514 -3814 186134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 221514 -3814 222134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 257514 460000 258134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 293514 460000 294134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 329514 460000 330134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 365514 460000 366134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 401514 460000 402134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 437514 -3814 438134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 473514 -3814 474134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 509514 -3814 510134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 545514 -3814 546134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 581514 -3814 582134 707750 4 vccd2
port 533 nsew
rlabel metal5 s -5846 -4774 589770 -4154 4 vdda1
port 534 nsew
rlabel metal5 s -6806 10306 590730 10926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 46306 590730 46926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 82306 590730 82926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 118306 590730 118926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 154306 590730 154926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 190306 590730 190926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 226306 590730 226926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 262306 590730 262926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 298306 590730 298926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 334306 590730 334926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 370306 590730 370926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 406306 590730 406926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 442306 590730 442926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 478306 590730 478926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 514306 590730 514926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 550306 590730 550926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 586306 590730 586926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 622306 590730 622926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 658306 590730 658926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 694306 590730 694926 4 vdda1
port 534 nsew
rlabel metal5 s -5846 708090 589770 708710 4 vdda1
port 534 nsew
rlabel metal4 s 261234 -5734 261854 336000 4 vdda1
port 534 nsew
rlabel metal4 s 297234 -5734 297854 336000 4 vdda1
port 534 nsew
rlabel metal4 s 333234 -5734 333854 336000 4 vdda1
port 534 nsew
rlabel metal4 s 369234 -5734 369854 336000 4 vdda1
port 534 nsew
rlabel metal4 s 405234 -5734 405854 336000 4 vdda1
port 534 nsew
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 534 nsew
rlabel metal4 s 589150 -4774 589770 708710 4 vdda1
port 534 nsew
rlabel metal4 s 9234 -5734 9854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 45234 -5734 45854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 81234 -5734 81854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 117234 -5734 117854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 153234 -5734 153854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 189234 -5734 189854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 225234 -5734 225854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 261234 460000 261854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 297234 460000 297854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 333234 460000 333854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 369234 460000 369854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 405234 460000 405854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 441234 -5734 441854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 477234 -5734 477854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 513234 -5734 513854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 549234 -5734 549854 709670 4 vdda1
port 534 nsew
rlabel metal5 s -7766 -6694 591690 -6074 4 vdda2
port 535 nsew
rlabel metal5 s -8726 14026 592650 14646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 50026 592650 50646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 86026 592650 86646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 122026 592650 122646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 158026 592650 158646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 194026 592650 194646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 230026 592650 230646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 266026 592650 266646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 302026 592650 302646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 338026 592650 338646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 374026 592650 374646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 410026 592650 410646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 446026 592650 446646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 482026 592650 482646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 518026 592650 518646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 554026 592650 554646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 590026 592650 590646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 626026 592650 626646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 662026 592650 662646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 698026 592650 698646 4 vdda2
port 535 nsew
rlabel metal5 s -7766 710010 591690 710630 4 vdda2
port 535 nsew
rlabel metal4 s 264954 -7654 265574 336000 4 vdda2
port 535 nsew
rlabel metal4 s 300954 -7654 301574 336000 4 vdda2
port 535 nsew
rlabel metal4 s 336954 -7654 337574 336000 4 vdda2
port 535 nsew
rlabel metal4 s 372954 -7654 373574 336000 4 vdda2
port 535 nsew
rlabel metal4 s 408954 -7654 409574 336000 4 vdda2
port 535 nsew
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 535 nsew
rlabel metal4 s 591070 -6694 591690 710630 4 vdda2
port 535 nsew
rlabel metal4 s 12954 -7654 13574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 48954 -7654 49574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 84954 -7654 85574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 120954 -7654 121574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 156954 -7654 157574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 192954 -7654 193574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 228954 -7654 229574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 264954 460000 265574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 300954 460000 301574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 336954 460000 337574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 372954 460000 373574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 408954 460000 409574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 444954 -7654 445574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 480954 -7654 481574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 516954 -7654 517574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 552954 -7654 553574 711590 4 vdda2
port 535 nsew
rlabel metal5 s -6806 -5734 590730 -5114 4 vssa1
port 536 nsew
rlabel metal5 s -6806 28306 590730 28926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 64306 590730 64926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 100306 590730 100926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 136306 590730 136926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 172306 590730 172926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 208306 590730 208926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 244306 590730 244926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 280306 590730 280926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 316306 590730 316926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 352306 590730 352926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 388306 590730 388926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 424306 590730 424926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 460306 590730 460926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 496306 590730 496926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 532306 590730 532926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 568306 590730 568926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 604306 590730 604926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 640306 590730 640926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 676306 590730 676926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 709050 590730 709670 4 vssa1
port 536 nsew
rlabel metal4 s 243234 -5734 243854 336000 4 vssa1
port 536 nsew
rlabel metal4 s 279234 -5734 279854 336000 4 vssa1
port 536 nsew
rlabel metal4 s 315234 -5734 315854 336000 4 vssa1
port 536 nsew
rlabel metal4 s 351234 -5734 351854 336000 4 vssa1
port 536 nsew
rlabel metal4 s 387234 -5734 387854 336000 4 vssa1
port 536 nsew
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 536 nsew
rlabel metal4 s 27234 -5734 27854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 63234 -5734 63854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 99234 -5734 99854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 135234 -5734 135854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 171234 -5734 171854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 207234 -5734 207854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 243234 460000 243854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 279234 460000 279854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 315234 460000 315854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 351234 460000 351854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 387234 460000 387854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 423234 -5734 423854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 459234 -5734 459854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 495234 -5734 495854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 531234 -5734 531854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 567234 -5734 567854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 590110 -5734 590730 709670 4 vssa1
port 536 nsew
rlabel metal5 s -8726 -7654 592650 -7034 4 vssa2
port 537 nsew
rlabel metal5 s -8726 32026 592650 32646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 68026 592650 68646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 104026 592650 104646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 140026 592650 140646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 176026 592650 176646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 212026 592650 212646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 248026 592650 248646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 284026 592650 284646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 320026 592650 320646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 356026 592650 356646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 392026 592650 392646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 428026 592650 428646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 464026 592650 464646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 500026 592650 500646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 536026 592650 536646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 572026 592650 572646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 608026 592650 608646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 644026 592650 644646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 680026 592650 680646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 710970 592650 711590 4 vssa2
port 537 nsew
rlabel metal4 s 246954 -7654 247574 336000 4 vssa2
port 537 nsew
rlabel metal4 s 282954 -7654 283574 336000 4 vssa2
port 537 nsew
rlabel metal4 s 318954 -7654 319574 336000 4 vssa2
port 537 nsew
rlabel metal4 s 354954 -7654 355574 336000 4 vssa2
port 537 nsew
rlabel metal4 s 390954 -7654 391574 336000 4 vssa2
port 537 nsew
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 537 nsew
rlabel metal4 s 30954 -7654 31574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 66954 -7654 67574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 102954 -7654 103574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 138954 -7654 139574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 174954 -7654 175574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 210954 -7654 211574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 246954 460000 247574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 282954 460000 283574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 318954 460000 319574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 354954 460000 355574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 390954 460000 391574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 426954 -7654 427574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 462954 -7654 463574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 498954 -7654 499574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 534954 -7654 535574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 570954 -7654 571574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 592030 -7654 592650 711590 4 vssa2
port 537 nsew
rlabel metal5 s -2966 -1894 586890 -1274 4 vssd1
port 538 nsew
rlabel metal5 s -2966 20866 586890 21486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 56866 586890 57486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 92866 586890 93486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 128866 586890 129486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 164866 586890 165486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 200866 586890 201486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 236866 586890 237486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 272866 586890 273486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 308866 586890 309486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 344866 586890 345486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 380866 586890 381486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 416866 586890 417486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 452866 586890 453486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 488866 586890 489486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 524866 586890 525486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 560866 586890 561486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 596866 586890 597486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 632866 586890 633486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 668866 586890 669486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 705210 586890 705830 4 vssd1
port 538 nsew
rlabel metal4 s 235794 -1894 236414 338000 4 vssd1
port 538 nsew
rlabel metal4 s 271794 -1894 272414 338000 4 vssd1
port 538 nsew
rlabel metal4 s 307794 -1894 308414 338000 4 vssd1
port 538 nsew
rlabel metal4 s 343794 -1894 344414 338000 4 vssd1
port 538 nsew
rlabel metal4 s 379794 -1894 380414 338000 4 vssd1
port 538 nsew
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 538 nsew
rlabel metal4 s 19794 -1894 20414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 55794 -1894 56414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 91794 -1894 92414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 127794 -1894 128414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 163794 -1894 164414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 199794 -1894 200414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 235794 458000 236414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 271794 458000 272414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 307794 458000 308414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 343794 458000 344414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 379794 458000 380414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 415794 -1894 416414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 451794 -1894 452414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 487794 -1894 488414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 523794 -1894 524414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 559794 -1894 560414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 586270 -1894 586890 705830 4 vssd1
port 538 nsew
rlabel metal5 s -4886 -3814 588810 -3194 4 vssd2
port 539 nsew
rlabel metal5 s -4886 24586 588810 25206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 60586 588810 61206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 96586 588810 97206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 132586 588810 133206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 168586 588810 169206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 204586 588810 205206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 240586 588810 241206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 276586 588810 277206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 312586 588810 313206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 348586 588810 349206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 384586 588810 385206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 420586 588810 421206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 456586 588810 457206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 492586 588810 493206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 528586 588810 529206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 564586 588810 565206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 600586 588810 601206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 636586 588810 637206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 672586 588810 673206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 707130 588810 707750 4 vssd2
port 539 nsew
rlabel metal4 s 239514 -3814 240134 336000 4 vssd2
port 539 nsew
rlabel metal4 s 275514 -3814 276134 336000 4 vssd2
port 539 nsew
rlabel metal4 s 311514 -3814 312134 336000 4 vssd2
port 539 nsew
rlabel metal4 s 347514 -3814 348134 336000 4 vssd2
port 539 nsew
rlabel metal4 s 383514 -3814 384134 336000 4 vssd2
port 539 nsew
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 539 nsew
rlabel metal4 s 23514 -3814 24134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 59514 -3814 60134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 95514 -3814 96134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 131514 -3814 132134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 167514 -3814 168134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 203514 -3814 204134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 239514 460000 240134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 275514 460000 276134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 311514 460000 312134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 347514 460000 348134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 383514 460000 384134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 419514 -3814 420134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 455514 -3814 456134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 491514 -3814 492134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 527514 -3814 528134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 563514 -3814 564134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 588190 -3814 588810 707750 4 vssd2
port 539 nsew
rlabel metal2 s 542 -960 654 480 4 wb_clk_i
port 540 nsew
rlabel metal2 s 1646 -960 1758 480 4 wb_rst_i
port 541 nsew
rlabel metal2 s 2842 -960 2954 480 4 wbs_ack_o
port 542 nsew
rlabel metal2 s 7626 -960 7738 480 4 wbs_adr_i[0]
port 543 nsew
rlabel metal2 s 47830 -960 47942 480 4 wbs_adr_i[10]
port 544 nsew
rlabel metal2 s 51326 -960 51438 480 4 wbs_adr_i[11]
port 545 nsew
rlabel metal2 s 54914 -960 55026 480 4 wbs_adr_i[12]
port 546 nsew
rlabel metal2 s 58410 -960 58522 480 4 wbs_adr_i[13]
port 547 nsew
rlabel metal2 s 61998 -960 62110 480 4 wbs_adr_i[14]
port 548 nsew
rlabel metal2 s 65494 -960 65606 480 4 wbs_adr_i[15]
port 549 nsew
rlabel metal2 s 69082 -960 69194 480 4 wbs_adr_i[16]
port 550 nsew
rlabel metal2 s 72578 -960 72690 480 4 wbs_adr_i[17]
port 551 nsew
rlabel metal2 s 76166 -960 76278 480 4 wbs_adr_i[18]
port 552 nsew
rlabel metal2 s 79662 -960 79774 480 4 wbs_adr_i[19]
port 553 nsew
rlabel metal2 s 12318 -960 12430 480 4 wbs_adr_i[1]
port 554 nsew
rlabel metal2 s 83250 -960 83362 480 4 wbs_adr_i[20]
port 555 nsew
rlabel metal2 s 86838 -960 86950 480 4 wbs_adr_i[21]
port 556 nsew
rlabel metal2 s 90334 -960 90446 480 4 wbs_adr_i[22]
port 557 nsew
rlabel metal2 s 93922 -960 94034 480 4 wbs_adr_i[23]
port 558 nsew
rlabel metal2 s 97418 -960 97530 480 4 wbs_adr_i[24]
port 559 nsew
rlabel metal2 s 101006 -960 101118 480 4 wbs_adr_i[25]
port 560 nsew
rlabel metal2 s 104502 -960 104614 480 4 wbs_adr_i[26]
port 561 nsew
rlabel metal2 s 108090 -960 108202 480 4 wbs_adr_i[27]
port 562 nsew
rlabel metal2 s 111586 -960 111698 480 4 wbs_adr_i[28]
port 563 nsew
rlabel metal2 s 115174 -960 115286 480 4 wbs_adr_i[29]
port 564 nsew
rlabel metal2 s 17010 -960 17122 480 4 wbs_adr_i[2]
port 565 nsew
rlabel metal2 s 118762 -960 118874 480 4 wbs_adr_i[30]
port 566 nsew
rlabel metal2 s 122258 -960 122370 480 4 wbs_adr_i[31]
port 567 nsew
rlabel metal2 s 21794 -960 21906 480 4 wbs_adr_i[3]
port 568 nsew
rlabel metal2 s 26486 -960 26598 480 4 wbs_adr_i[4]
port 569 nsew
rlabel metal2 s 30074 -960 30186 480 4 wbs_adr_i[5]
port 570 nsew
rlabel metal2 s 33570 -960 33682 480 4 wbs_adr_i[6]
port 571 nsew
rlabel metal2 s 37158 -960 37270 480 4 wbs_adr_i[7]
port 572 nsew
rlabel metal2 s 40654 -960 40766 480 4 wbs_adr_i[8]
port 573 nsew
rlabel metal2 s 44242 -960 44354 480 4 wbs_adr_i[9]
port 574 nsew
rlabel metal2 s 4038 -960 4150 480 4 wbs_cyc_i
port 575 nsew
rlabel metal2 s 8730 -960 8842 480 4 wbs_dat_i[0]
port 576 nsew
rlabel metal2 s 48934 -960 49046 480 4 wbs_dat_i[10]
port 577 nsew
rlabel metal2 s 52522 -960 52634 480 4 wbs_dat_i[11]
port 578 nsew
rlabel metal2 s 56018 -960 56130 480 4 wbs_dat_i[12]
port 579 nsew
rlabel metal2 s 59606 -960 59718 480 4 wbs_dat_i[13]
port 580 nsew
rlabel metal2 s 63194 -960 63306 480 4 wbs_dat_i[14]
port 581 nsew
rlabel metal2 s 66690 -960 66802 480 4 wbs_dat_i[15]
port 582 nsew
rlabel metal2 s 70278 -960 70390 480 4 wbs_dat_i[16]
port 583 nsew
rlabel metal2 s 73774 -960 73886 480 4 wbs_dat_i[17]
port 584 nsew
rlabel metal2 s 77362 -960 77474 480 4 wbs_dat_i[18]
port 585 nsew
rlabel metal2 s 80858 -960 80970 480 4 wbs_dat_i[19]
port 586 nsew
rlabel metal2 s 13514 -960 13626 480 4 wbs_dat_i[1]
port 587 nsew
rlabel metal2 s 84446 -960 84558 480 4 wbs_dat_i[20]
port 588 nsew
rlabel metal2 s 87942 -960 88054 480 4 wbs_dat_i[21]
port 589 nsew
rlabel metal2 s 91530 -960 91642 480 4 wbs_dat_i[22]
port 590 nsew
rlabel metal2 s 95118 -960 95230 480 4 wbs_dat_i[23]
port 591 nsew
rlabel metal2 s 98614 -960 98726 480 4 wbs_dat_i[24]
port 592 nsew
rlabel metal2 s 102202 -960 102314 480 4 wbs_dat_i[25]
port 593 nsew
rlabel metal2 s 105698 -960 105810 480 4 wbs_dat_i[26]
port 594 nsew
rlabel metal2 s 109286 -960 109398 480 4 wbs_dat_i[27]
port 595 nsew
rlabel metal2 s 112782 -960 112894 480 4 wbs_dat_i[28]
port 596 nsew
rlabel metal2 s 116370 -960 116482 480 4 wbs_dat_i[29]
port 597 nsew
rlabel metal2 s 18206 -960 18318 480 4 wbs_dat_i[2]
port 598 nsew
rlabel metal2 s 119866 -960 119978 480 4 wbs_dat_i[30]
port 599 nsew
rlabel metal2 s 123454 -960 123566 480 4 wbs_dat_i[31]
port 600 nsew
rlabel metal2 s 22990 -960 23102 480 4 wbs_dat_i[3]
port 601 nsew
rlabel metal2 s 27682 -960 27794 480 4 wbs_dat_i[4]
port 602 nsew
rlabel metal2 s 31270 -960 31382 480 4 wbs_dat_i[5]
port 603 nsew
rlabel metal2 s 34766 -960 34878 480 4 wbs_dat_i[6]
port 604 nsew
rlabel metal2 s 38354 -960 38466 480 4 wbs_dat_i[7]
port 605 nsew
rlabel metal2 s 41850 -960 41962 480 4 wbs_dat_i[8]
port 606 nsew
rlabel metal2 s 45438 -960 45550 480 4 wbs_dat_i[9]
port 607 nsew
rlabel metal2 s 9926 -960 10038 480 4 wbs_dat_o[0]
port 608 nsew
rlabel metal2 s 50130 -960 50242 480 4 wbs_dat_o[10]
port 609 nsew
rlabel metal2 s 53718 -960 53830 480 4 wbs_dat_o[11]
port 610 nsew
rlabel metal2 s 57214 -960 57326 480 4 wbs_dat_o[12]
port 611 nsew
rlabel metal2 s 60802 -960 60914 480 4 wbs_dat_o[13]
port 612 nsew
rlabel metal2 s 64298 -960 64410 480 4 wbs_dat_o[14]
port 613 nsew
rlabel metal2 s 67886 -960 67998 480 4 wbs_dat_o[15]
port 614 nsew
rlabel metal2 s 71474 -960 71586 480 4 wbs_dat_o[16]
port 615 nsew
rlabel metal2 s 74970 -960 75082 480 4 wbs_dat_o[17]
port 616 nsew
rlabel metal2 s 78558 -960 78670 480 4 wbs_dat_o[18]
port 617 nsew
rlabel metal2 s 82054 -960 82166 480 4 wbs_dat_o[19]
port 618 nsew
rlabel metal2 s 14710 -960 14822 480 4 wbs_dat_o[1]
port 619 nsew
rlabel metal2 s 85642 -960 85754 480 4 wbs_dat_o[20]
port 620 nsew
rlabel metal2 s 89138 -960 89250 480 4 wbs_dat_o[21]
port 621 nsew
rlabel metal2 s 92726 -960 92838 480 4 wbs_dat_o[22]
port 622 nsew
rlabel metal2 s 96222 -960 96334 480 4 wbs_dat_o[23]
port 623 nsew
rlabel metal2 s 99810 -960 99922 480 4 wbs_dat_o[24]
port 624 nsew
rlabel metal2 s 103306 -960 103418 480 4 wbs_dat_o[25]
port 625 nsew
rlabel metal2 s 106894 -960 107006 480 4 wbs_dat_o[26]
port 626 nsew
rlabel metal2 s 110482 -960 110594 480 4 wbs_dat_o[27]
port 627 nsew
rlabel metal2 s 113978 -960 114090 480 4 wbs_dat_o[28]
port 628 nsew
rlabel metal2 s 117566 -960 117678 480 4 wbs_dat_o[29]
port 629 nsew
rlabel metal2 s 19402 -960 19514 480 4 wbs_dat_o[2]
port 630 nsew
rlabel metal2 s 121062 -960 121174 480 4 wbs_dat_o[30]
port 631 nsew
rlabel metal2 s 124650 -960 124762 480 4 wbs_dat_o[31]
port 632 nsew
rlabel metal2 s 24186 -960 24298 480 4 wbs_dat_o[3]
port 633 nsew
rlabel metal2 s 28878 -960 28990 480 4 wbs_dat_o[4]
port 634 nsew
rlabel metal2 s 32374 -960 32486 480 4 wbs_dat_o[5]
port 635 nsew
rlabel metal2 s 35962 -960 36074 480 4 wbs_dat_o[6]
port 636 nsew
rlabel metal2 s 39550 -960 39662 480 4 wbs_dat_o[7]
port 637 nsew
rlabel metal2 s 43046 -960 43158 480 4 wbs_dat_o[8]
port 638 nsew
rlabel metal2 s 46634 -960 46746 480 4 wbs_dat_o[9]
port 639 nsew
rlabel metal2 s 11122 -960 11234 480 4 wbs_sel_i[0]
port 640 nsew
rlabel metal2 s 15906 -960 16018 480 4 wbs_sel_i[1]
port 641 nsew
rlabel metal2 s 20598 -960 20710 480 4 wbs_sel_i[2]
port 642 nsew
rlabel metal2 s 25290 -960 25402 480 4 wbs_sel_i[3]
port 643 nsew
rlabel metal2 s 5234 -960 5346 480 4 wbs_stb_i
port 644 nsew
rlabel metal2 s 6430 -960 6542 480 4 wbs_we_i
port 645 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
