magic
tech sky130A
magscale 1 2
timestamp 1634570663
<< checkpaint >>
rect -12658 -11586 596582 715522
<< locali >>
rect 263275 379729 263517 379763
rect 253213 377791 253247 377893
rect 253121 377655 253155 377757
rect 238585 376771 238619 377553
rect 239229 376839 239263 377553
rect 240793 376975 240827 377553
rect 241621 376907 241655 377553
rect 247601 377247 247635 377553
rect 284861 377111 284895 377417
rect 288541 377043 288575 377349
rect 290657 377179 290691 377349
rect 236561 337603 236595 337977
rect 239413 335359 239447 336617
rect 236009 331415 236043 332061
rect 230305 330191 230339 330565
rect 245025 329647 245059 337773
rect 249165 336379 249199 336413
rect 249015 336345 249199 336379
rect 249107 336209 249199 336243
rect 248797 335359 248831 335869
rect 248981 335835 249015 336141
rect 249165 336039 249199 336209
rect 249257 336107 249291 336277
rect 249073 335903 249107 336005
rect 248889 335495 248923 335801
rect 248981 335665 249165 335699
rect 248981 335631 249015 335665
rect 251281 335427 251315 337841
rect 252017 336243 252051 336685
rect 248705 335019 248739 335325
rect 251373 335019 251407 335393
rect 255789 330327 255823 337773
rect 264069 335835 264103 337909
rect 264253 330871 264287 337909
rect 267565 331891 267599 337909
rect 270141 328695 270175 337841
rect 271337 334543 271371 337841
rect 271521 332979 271555 337841
rect 273453 337535 273487 337909
rect 274925 337535 274959 337841
rect 273913 336515 273947 336617
rect 272809 335767 272843 335937
rect 273085 335699 273119 336277
rect 273177 335903 273211 336209
rect 272993 335495 273027 335665
rect 273269 335495 273303 335733
rect 274005 335699 274039 336481
rect 276765 333183 276799 337909
rect 278053 336175 278087 336345
rect 278145 335563 278179 335937
rect 278237 333931 278271 337841
rect 278605 336175 278639 337909
rect 280077 336243 280111 337977
rect 280445 337195 280479 337909
rect 283665 336991 283699 337909
rect 282561 336685 282871 336719
rect 280169 335495 280203 335801
rect 281365 335223 281399 335665
rect 282377 333115 282411 336277
rect 282469 335495 282503 336413
rect 282561 335835 282595 336685
rect 282469 335461 282653 335495
rect 282745 335427 282779 336617
rect 282837 336311 282871 336685
rect 283205 335767 283239 336413
rect 283113 335359 283147 335665
rect 283297 335563 283331 335733
rect 284033 332503 284067 337909
rect 284401 334611 284435 337773
rect 285505 335223 285539 335733
rect 286057 334883 286091 337773
rect 287713 337195 287747 337841
rect 289277 336107 289311 336413
rect 289369 336107 289403 337773
rect 286333 335427 286367 335665
rect 288541 335563 288575 335937
rect 292405 335495 292439 335665
rect 292221 335223 292255 335325
rect 292497 335223 292531 336685
rect 292589 335563 292623 336685
rect 292681 335223 292715 335529
rect 294061 335359 294095 335597
rect 294153 335427 294187 335597
rect 289921 334985 290013 335019
rect 289921 334611 289955 334985
rect 294245 329103 294279 337841
rect 294337 332027 294371 337909
rect 294797 335971 294831 336481
rect 294889 336039 294923 336481
rect 294797 335937 295383 335971
rect 294555 335869 295257 335903
rect 295349 335563 295383 335937
rect 294831 335529 295015 335563
rect 294981 335427 295015 335529
rect 297373 335495 297407 336005
rect 294739 335325 295257 335359
rect 295073 334815 295107 335257
rect 234997 323595 235031 326689
rect 235825 326587 235859 326689
rect 290657 326655 290691 326757
rect 280629 326315 280663 326553
rect 582389 46359 582423 378165
rect 582481 73015 582515 378233
rect 582573 86207 582607 376737
rect 582665 99535 582699 378369
rect 582757 112863 582791 376805
rect 582849 126055 582883 378301
rect 232053 4811 232087 4913
rect 88901 3995 88935 4097
rect 233341 3757 233985 3791
rect 233341 3587 233375 3757
rect 102241 3043 102275 3281
rect 102333 2907 102367 3145
rect 128921 2941 129105 2975
rect 128921 2839 128955 2941
rect 229293 2839 229327 3417
rect 436845 3315 436879 4029
rect 456073 3859 456107 3961
rect 452393 3383 452427 3757
rect 582941 3247 582975 336753
rect 583033 152711 583067 376941
rect 583125 165903 583159 376873
rect 409245 3009 409521 3043
rect 409245 2975 409279 3009
<< viali >>
rect 263241 379729 263275 379763
rect 263517 379729 263551 379763
rect 582665 378369 582699 378403
rect 582481 378233 582515 378267
rect 582389 378165 582423 378199
rect 253213 377893 253247 377927
rect 253121 377757 253155 377791
rect 253213 377757 253247 377791
rect 253121 377621 253155 377655
rect 238585 377553 238619 377587
rect 239229 377553 239263 377587
rect 240793 377553 240827 377587
rect 240793 376941 240827 376975
rect 241621 377553 241655 377587
rect 247601 377553 247635 377587
rect 247601 377213 247635 377247
rect 284861 377417 284895 377451
rect 284861 377077 284895 377111
rect 288541 377349 288575 377383
rect 290657 377349 290691 377383
rect 290657 377145 290691 377179
rect 288541 377009 288575 377043
rect 241621 376873 241655 376907
rect 239229 376805 239263 376839
rect 238585 376737 238619 376771
rect 236561 337977 236595 338011
rect 280077 337977 280111 338011
rect 264069 337909 264103 337943
rect 251281 337841 251315 337875
rect 236561 337569 236595 337603
rect 245025 337773 245059 337807
rect 239413 336617 239447 336651
rect 239413 335325 239447 335359
rect 236009 332061 236043 332095
rect 236009 331381 236043 331415
rect 230305 330565 230339 330599
rect 230305 330157 230339 330191
rect 249165 336413 249199 336447
rect 248981 336345 249015 336379
rect 249257 336277 249291 336311
rect 249073 336209 249107 336243
rect 248981 336141 249015 336175
rect 248797 335869 248831 335903
rect 249257 336073 249291 336107
rect 249073 336005 249107 336039
rect 249165 336005 249199 336039
rect 249073 335869 249107 335903
rect 248889 335801 248923 335835
rect 248981 335801 249015 335835
rect 249165 335665 249199 335699
rect 248981 335597 249015 335631
rect 248889 335461 248923 335495
rect 255789 337773 255823 337807
rect 252017 336685 252051 336719
rect 252017 336209 252051 336243
rect 251281 335393 251315 335427
rect 251373 335393 251407 335427
rect 248705 335325 248739 335359
rect 248797 335325 248831 335359
rect 248705 334985 248739 335019
rect 251373 334985 251407 335019
rect 264069 335801 264103 335835
rect 264253 337909 264287 337943
rect 267565 337909 267599 337943
rect 273453 337909 273487 337943
rect 267565 331857 267599 331891
rect 270141 337841 270175 337875
rect 264253 330837 264287 330871
rect 255789 330293 255823 330327
rect 245025 329613 245059 329647
rect 271337 337841 271371 337875
rect 271337 334509 271371 334543
rect 271521 337841 271555 337875
rect 276765 337909 276799 337943
rect 273453 337501 273487 337535
rect 274925 337841 274959 337875
rect 274925 337501 274959 337535
rect 273913 336617 273947 336651
rect 273913 336481 273947 336515
rect 274005 336481 274039 336515
rect 273085 336277 273119 336311
rect 272809 335937 272843 335971
rect 272809 335733 272843 335767
rect 273177 336209 273211 336243
rect 273177 335869 273211 335903
rect 272993 335665 273027 335699
rect 273085 335665 273119 335699
rect 273269 335733 273303 335767
rect 272993 335461 273027 335495
rect 274005 335665 274039 335699
rect 273269 335461 273303 335495
rect 278605 337909 278639 337943
rect 278237 337841 278271 337875
rect 278053 336345 278087 336379
rect 278053 336141 278087 336175
rect 278145 335937 278179 335971
rect 278145 335529 278179 335563
rect 280445 337909 280479 337943
rect 280445 337161 280479 337195
rect 283665 337909 283699 337943
rect 283665 336957 283699 336991
rect 284033 337909 284067 337943
rect 282469 336413 282503 336447
rect 280077 336209 280111 336243
rect 282377 336277 282411 336311
rect 278605 336141 278639 336175
rect 280169 335801 280203 335835
rect 280169 335461 280203 335495
rect 281365 335665 281399 335699
rect 281365 335189 281399 335223
rect 278237 333897 278271 333931
rect 276765 333149 276799 333183
rect 282561 335801 282595 335835
rect 282745 336617 282779 336651
rect 282653 335461 282687 335495
rect 282837 336277 282871 336311
rect 283205 336413 283239 336447
rect 283205 335733 283239 335767
rect 283297 335733 283331 335767
rect 282745 335393 282779 335427
rect 283113 335665 283147 335699
rect 283297 335529 283331 335563
rect 283113 335325 283147 335359
rect 282377 333081 282411 333115
rect 271521 332945 271555 332979
rect 294337 337909 294371 337943
rect 287713 337841 287747 337875
rect 284401 337773 284435 337807
rect 286057 337773 286091 337807
rect 285505 335733 285539 335767
rect 285505 335189 285539 335223
rect 294245 337841 294279 337875
rect 287713 337161 287747 337195
rect 289369 337773 289403 337807
rect 289277 336413 289311 336447
rect 289277 336073 289311 336107
rect 289369 336073 289403 336107
rect 292497 336685 292531 336719
rect 288541 335937 288575 335971
rect 286333 335665 286367 335699
rect 288541 335529 288575 335563
rect 292405 335665 292439 335699
rect 292405 335461 292439 335495
rect 286333 335393 286367 335427
rect 292221 335325 292255 335359
rect 292221 335189 292255 335223
rect 292589 336685 292623 336719
rect 294061 335597 294095 335631
rect 292589 335529 292623 335563
rect 292681 335529 292715 335563
rect 292497 335189 292531 335223
rect 294153 335597 294187 335631
rect 294153 335393 294187 335427
rect 294061 335325 294095 335359
rect 292681 335189 292715 335223
rect 286057 334849 286091 334883
rect 290013 334985 290047 335019
rect 284401 334577 284435 334611
rect 289921 334577 289955 334611
rect 284033 332469 284067 332503
rect 294797 336481 294831 336515
rect 294889 336481 294923 336515
rect 294889 336005 294923 336039
rect 297373 336005 297407 336039
rect 294521 335869 294555 335903
rect 295257 335869 295291 335903
rect 294797 335529 294831 335563
rect 295349 335529 295383 335563
rect 297373 335461 297407 335495
rect 294981 335393 295015 335427
rect 294705 335325 294739 335359
rect 295257 335325 295291 335359
rect 295073 335257 295107 335291
rect 295073 334781 295107 334815
rect 294337 331993 294371 332027
rect 294245 329069 294279 329103
rect 270141 328661 270175 328695
rect 290657 326757 290691 326791
rect 234997 326689 235031 326723
rect 235825 326689 235859 326723
rect 290657 326621 290691 326655
rect 235825 326553 235859 326587
rect 280629 326553 280663 326587
rect 280629 326281 280663 326315
rect 234997 323561 235031 323595
rect 582573 376737 582607 376771
rect 582849 378301 582883 378335
rect 582757 376805 582791 376839
rect 583033 376941 583067 376975
rect 582849 126021 582883 126055
rect 582941 336753 582975 336787
rect 582757 112829 582791 112863
rect 582665 99501 582699 99535
rect 582573 86173 582607 86207
rect 582481 72981 582515 73015
rect 582389 46325 582423 46359
rect 232053 4913 232087 4947
rect 232053 4777 232087 4811
rect 88901 4097 88935 4131
rect 88901 3961 88935 3995
rect 436845 4029 436879 4063
rect 233985 3757 234019 3791
rect 233341 3553 233375 3587
rect 229293 3417 229327 3451
rect 102241 3281 102275 3315
rect 102241 3009 102275 3043
rect 102333 3145 102367 3179
rect 102333 2873 102367 2907
rect 129105 2941 129139 2975
rect 128921 2805 128955 2839
rect 456073 3961 456107 3995
rect 456073 3825 456107 3859
rect 452393 3757 452427 3791
rect 452393 3349 452427 3383
rect 436845 3281 436879 3315
rect 583125 376873 583159 376907
rect 583125 165869 583159 165903
rect 583033 152677 583067 152711
rect 582941 3213 582975 3247
rect 409521 3009 409555 3043
rect 409245 2941 409279 2975
rect 229293 2805 229327 2839
<< metal1 >>
rect 263318 700952 263324 701004
rect 263376 700992 263382 701004
rect 397454 700992 397460 701004
rect 263376 700964 397460 700992
rect 263376 700952 263382 700964
rect 397454 700952 397460 700964
rect 397512 700952 397518 701004
rect 263502 700884 263508 700936
rect 263560 700924 263566 700936
rect 413646 700924 413652 700936
rect 263560 700896 413652 700924
rect 263560 700884 263566 700896
rect 413646 700884 413652 700896
rect 413704 700884 413710 700936
rect 262030 700816 262036 700868
rect 262088 700856 262094 700868
rect 429838 700856 429844 700868
rect 262088 700828 429844 700856
rect 262088 700816 262094 700828
rect 429838 700816 429844 700828
rect 429896 700816 429902 700868
rect 72970 700748 72976 700800
rect 73028 700788 73034 700800
rect 269482 700788 269488 700800
rect 73028 700760 269488 700788
rect 73028 700748 73034 700760
rect 269482 700748 269488 700760
rect 269540 700748 269546 700800
rect 262122 700680 262128 700732
rect 262180 700720 262186 700732
rect 462314 700720 462320 700732
rect 262180 700692 462320 700720
rect 262180 700680 262186 700692
rect 462314 700680 462320 700692
rect 462372 700680 462378 700732
rect 261938 700612 261944 700664
rect 261996 700652 262002 700664
rect 478506 700652 478512 700664
rect 261996 700624 478512 700652
rect 261996 700612 262002 700624
rect 478506 700612 478512 700624
rect 478564 700612 478570 700664
rect 260650 700544 260656 700596
rect 260708 700584 260714 700596
rect 494790 700584 494796 700596
rect 260708 700556 494796 700584
rect 260708 700544 260714 700556
rect 494790 700544 494796 700556
rect 494848 700544 494854 700596
rect 8110 700476 8116 700528
rect 8168 700516 8174 700528
rect 271874 700516 271880 700528
rect 8168 700488 271880 700516
rect 8168 700476 8174 700488
rect 271874 700476 271880 700488
rect 271932 700476 271938 700528
rect 259362 700408 259368 700460
rect 259420 700448 259426 700460
rect 527174 700448 527180 700460
rect 259420 700420 527180 700448
rect 259420 700408 259426 700420
rect 527174 700408 527180 700420
rect 527232 700408 527238 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 41322 700380 41328 700392
rect 40552 700352 41328 700380
rect 40552 700340 40558 700352
rect 41322 700340 41328 700352
rect 41380 700340 41386 700392
rect 260742 700340 260748 700392
rect 260800 700380 260806 700392
rect 543458 700380 543464 700392
rect 260800 700352 543464 700380
rect 260800 700340 260806 700352
rect 543458 700340 543464 700352
rect 543516 700340 543522 700392
rect 259270 700272 259276 700324
rect 259328 700312 259334 700324
rect 559650 700312 559656 700324
rect 259328 700284 559656 700312
rect 259328 700272 259334 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 137830 700204 137836 700256
rect 137888 700244 137894 700256
rect 267918 700244 267924 700256
rect 137888 700216 267924 700244
rect 137888 700204 137894 700216
rect 267918 700204 267924 700216
rect 267976 700204 267982 700256
rect 263410 700136 263416 700188
rect 263468 700176 263474 700188
rect 364978 700176 364984 700188
rect 263468 700148 364984 700176
rect 263468 700136 263474 700148
rect 364978 700136 364984 700148
rect 365036 700136 365042 700188
rect 264790 700068 264796 700120
rect 264848 700108 264854 700120
rect 348786 700108 348792 700120
rect 264848 700080 348792 700108
rect 264848 700068 264854 700080
rect 348786 700068 348792 700080
rect 348844 700068 348850 700120
rect 264882 700000 264888 700052
rect 264940 700040 264946 700052
rect 332502 700040 332508 700052
rect 264940 700012 332508 700040
rect 264940 700000 264946 700012
rect 332502 700000 332508 700012
rect 332560 700000 332566 700052
rect 202782 699932 202788 699984
rect 202840 699972 202846 699984
rect 266446 699972 266452 699984
rect 202840 699944 266452 699972
rect 202840 699932 202846 699944
rect 266446 699932 266452 699944
rect 266504 699932 266510 699984
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 170306 699660 170312 699712
rect 170364 699700 170370 699712
rect 171042 699700 171048 699712
rect 170364 699672 171048 699700
rect 170364 699660 170370 699672
rect 171042 699660 171048 699672
rect 171100 699660 171106 699712
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 235902 699700 235908 699712
rect 235224 699672 235908 699700
rect 235224 699660 235230 699672
rect 235902 699660 235908 699672
rect 235960 699660 235966 699712
rect 266262 699660 266268 699712
rect 266320 699700 266326 699712
rect 267642 699700 267648 699712
rect 266320 699672 267648 699700
rect 266320 699660 266326 699672
rect 267642 699660 267648 699672
rect 267700 699660 267706 699712
rect 257982 696940 257988 696992
rect 258040 696980 258046 696992
rect 580166 696980 580172 696992
rect 258040 696952 580172 696980
rect 258040 696940 258046 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 259178 683136 259184 683188
rect 259236 683176 259242 683188
rect 580166 683176 580172 683188
rect 259236 683148 580172 683176
rect 259236 683136 259242 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 257890 670692 257896 670744
rect 257948 670732 257954 670744
rect 580166 670732 580172 670744
rect 257948 670704 580172 670732
rect 257948 670692 257954 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3142 656888 3148 656940
rect 3200 656928 3206 656940
rect 273438 656928 273444 656940
rect 3200 656900 273444 656928
rect 3200 656888 3206 656900
rect 273438 656888 273444 656900
rect 273496 656888 273502 656940
rect 256602 643084 256608 643136
rect 256660 643124 256666 643136
rect 580166 643124 580172 643136
rect 256660 643096 580172 643124
rect 256660 643084 256666 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 257798 630640 257804 630692
rect 257856 630680 257862 630692
rect 580166 630680 580172 630692
rect 257856 630652 580172 630680
rect 257856 630640 257862 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 256510 616836 256516 616888
rect 256568 616876 256574 616888
rect 580166 616876 580172 616888
rect 256568 616848 580172 616876
rect 256568 616836 256574 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3326 605820 3332 605872
rect 3384 605860 3390 605872
rect 274726 605860 274732 605872
rect 3384 605832 274732 605860
rect 3384 605820 3390 605832
rect 274726 605820 274732 605832
rect 274784 605820 274790 605872
rect 255222 590656 255228 590708
rect 255280 590696 255286 590708
rect 579798 590696 579804 590708
rect 255280 590668 579804 590696
rect 255280 590656 255286 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 255130 576852 255136 576904
rect 255188 576892 255194 576904
rect 580166 576892 580172 576904
rect 255188 576864 580172 576892
rect 255188 576852 255194 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 255038 563048 255044 563100
rect 255096 563088 255102 563100
rect 579798 563088 579804 563100
rect 255096 563060 579804 563088
rect 255096 563048 255102 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3142 553392 3148 553444
rect 3200 553432 3206 553444
rect 276382 553432 276388 553444
rect 3200 553404 276388 553432
rect 3200 553392 3206 553404
rect 276382 553392 276388 553404
rect 276440 553392 276446 553444
rect 253842 536800 253848 536852
rect 253900 536840 253906 536852
rect 580166 536840 580172 536852
rect 253900 536812 580172 536840
rect 253900 536800 253906 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 253750 524424 253756 524476
rect 253808 524464 253814 524476
rect 580166 524464 580172 524476
rect 253808 524436 580172 524464
rect 253808 524424 253814 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 252462 510620 252468 510672
rect 252520 510660 252526 510672
rect 580166 510660 580172 510672
rect 252520 510632 580172 510660
rect 252520 510620 252526 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3234 500964 3240 501016
rect 3292 501004 3298 501016
rect 277486 501004 277492 501016
rect 3292 500976 277492 501004
rect 3292 500964 3298 500976
rect 277486 500964 277492 500976
rect 277544 500964 277550 501016
rect 252370 484372 252376 484424
rect 252428 484412 252434 484424
rect 580166 484412 580172 484424
rect 252428 484384 580172 484412
rect 252428 484372 252434 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 252278 470568 252284 470620
rect 252336 470608 252342 470620
rect 579982 470608 579988 470620
rect 252336 470580 579988 470608
rect 252336 470568 252342 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 251082 456764 251088 456816
rect 251140 456804 251146 456816
rect 580166 456804 580172 456816
rect 251140 456776 580172 456804
rect 251140 456764 251146 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 278958 448576 278964 448588
rect 3200 448548 278964 448576
rect 3200 448536 3206 448548
rect 278958 448536 278964 448548
rect 279016 448536 279022 448588
rect 250990 430584 250996 430636
rect 251048 430624 251054 430636
rect 580166 430624 580172 430636
rect 251048 430596 580172 430624
rect 251048 430584 251054 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 250898 418140 250904 418192
rect 250956 418180 250962 418192
rect 580166 418180 580172 418192
rect 250956 418152 580172 418180
rect 250956 418140 250962 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 249702 404336 249708 404388
rect 249760 404376 249766 404388
rect 580166 404376 580172 404388
rect 249760 404348 580172 404376
rect 249760 404336 249766 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 2958 397468 2964 397520
rect 3016 397508 3022 397520
rect 281074 397508 281080 397520
rect 3016 397480 281080 397508
rect 3016 397468 3022 397480
rect 281074 397468 281080 397480
rect 281132 397468 281138 397520
rect 3602 380808 3608 380860
rect 3660 380848 3666 380860
rect 274266 380848 274272 380860
rect 3660 380820 274272 380848
rect 3660 380808 3666 380820
rect 274266 380808 274272 380820
rect 274324 380808 274330 380860
rect 3510 380740 3516 380792
rect 3568 380780 3574 380792
rect 273806 380780 273812 380792
rect 3568 380752 273812 380780
rect 3568 380740 3574 380752
rect 273806 380740 273812 380752
rect 273864 380740 273870 380792
rect 3694 380672 3700 380724
rect 3752 380712 3758 380724
rect 275370 380712 275376 380724
rect 3752 380684 275376 380712
rect 3752 380672 3758 380684
rect 275370 380672 275376 380684
rect 275428 380672 275434 380724
rect 3878 380604 3884 380656
rect 3936 380644 3942 380656
rect 276934 380644 276940 380656
rect 3936 380616 276940 380644
rect 3936 380604 3942 380616
rect 276934 380604 276940 380616
rect 276992 380604 276998 380656
rect 3786 380536 3792 380588
rect 3844 380576 3850 380588
rect 276014 380576 276020 380588
rect 3844 380548 276020 380576
rect 3844 380536 3850 380548
rect 276014 380536 276020 380548
rect 276072 380536 276078 380588
rect 3970 380468 3976 380520
rect 4028 380508 4034 380520
rect 277578 380508 277584 380520
rect 4028 380480 277584 380508
rect 4028 380468 4034 380480
rect 277578 380468 277584 380480
rect 277636 380468 277642 380520
rect 4062 380400 4068 380452
rect 4120 380440 4126 380452
rect 278774 380440 278780 380452
rect 4120 380412 278780 380440
rect 4120 380400 4126 380412
rect 278774 380400 278780 380412
rect 278832 380400 278838 380452
rect 3326 380332 3332 380384
rect 3384 380372 3390 380384
rect 279050 380372 279056 380384
rect 3384 380344 279056 380372
rect 3384 380332 3390 380344
rect 279050 380332 279056 380344
rect 279108 380332 279114 380384
rect 3234 380264 3240 380316
rect 3292 380304 3298 380316
rect 280154 380304 280160 380316
rect 3292 380276 280160 380304
rect 3292 380264 3298 380276
rect 280154 380264 280160 380276
rect 280212 380264 280218 380316
rect 3142 380196 3148 380248
rect 3200 380236 3206 380248
rect 280614 380236 280620 380248
rect 3200 380208 280620 380236
rect 3200 380196 3206 380208
rect 280614 380196 280620 380208
rect 280672 380196 280678 380248
rect 3050 380128 3056 380180
rect 3108 380168 3114 380180
rect 281718 380168 281724 380180
rect 3108 380140 281724 380168
rect 3108 380128 3114 380140
rect 281718 380128 281724 380140
rect 281776 380128 281782 380180
rect 41322 380060 41328 380112
rect 41380 380100 41386 380112
rect 271138 380100 271144 380112
rect 41380 380072 271144 380100
rect 41380 380060 41386 380072
rect 271138 380060 271144 380072
rect 271196 380060 271202 380112
rect 106182 379992 106188 380044
rect 106240 380032 106246 380044
rect 269574 380032 269580 380044
rect 106240 380004 269580 380032
rect 106240 379992 106246 380004
rect 269574 379992 269580 380004
rect 269632 379992 269638 380044
rect 89622 379924 89628 379976
rect 89680 379964 89686 379976
rect 270586 379964 270592 379976
rect 89680 379936 270592 379964
rect 89680 379924 89686 379936
rect 270586 379924 270592 379936
rect 270644 379924 270650 379976
rect 154482 379856 154488 379908
rect 154540 379896 154546 379908
rect 269114 379896 269120 379908
rect 154540 379868 269120 379896
rect 154540 379856 154546 379868
rect 269114 379856 269120 379868
rect 269172 379856 269178 379908
rect 171042 379788 171048 379840
rect 171100 379828 171106 379840
rect 171100 379800 258580 379828
rect 171100 379788 171106 379800
rect 219342 379720 219348 379772
rect 219400 379760 219406 379772
rect 258552 379760 258580 379800
rect 258626 379788 258632 379840
rect 258684 379828 258690 379840
rect 259178 379828 259184 379840
rect 258684 379800 259184 379828
rect 258684 379788 258690 379800
rect 259178 379788 259184 379800
rect 259236 379788 259242 379840
rect 260190 379788 260196 379840
rect 260248 379828 260254 379840
rect 260742 379828 260748 379840
rect 260248 379800 260748 379828
rect 260248 379788 260254 379800
rect 260742 379788 260748 379800
rect 260800 379788 260806 379840
rect 261294 379788 261300 379840
rect 261352 379828 261358 379840
rect 262122 379828 262128 379840
rect 261352 379800 262128 379828
rect 261352 379788 261358 379800
rect 262122 379788 262128 379800
rect 262180 379788 262186 379840
rect 262858 379788 262864 379840
rect 262916 379828 262922 379840
rect 263318 379828 263324 379840
rect 262916 379800 263324 379828
rect 262916 379788 262922 379800
rect 263318 379788 263324 379800
rect 263376 379788 263382 379840
rect 267734 379828 267740 379840
rect 263428 379800 267740 379828
rect 263229 379763 263287 379769
rect 263229 379760 263241 379763
rect 219400 379732 258074 379760
rect 258552 379732 263241 379760
rect 219400 379720 219406 379732
rect 250254 379652 250260 379704
rect 250312 379692 250318 379704
rect 250990 379692 250996 379704
rect 250312 379664 250996 379692
rect 250312 379652 250318 379664
rect 250990 379652 250996 379664
rect 251048 379652 251054 379704
rect 251818 379652 251824 379704
rect 251876 379692 251882 379704
rect 252370 379692 252376 379704
rect 251876 379664 252376 379692
rect 251876 379652 251882 379664
rect 252370 379652 252376 379664
rect 252428 379652 252434 379704
rect 253382 379652 253388 379704
rect 253440 379692 253446 379704
rect 253842 379692 253848 379704
rect 253440 379664 253848 379692
rect 253440 379652 253446 379664
rect 253842 379652 253848 379664
rect 253900 379652 253906 379704
rect 254394 379652 254400 379704
rect 254452 379692 254458 379704
rect 255038 379692 255044 379704
rect 254452 379664 255044 379692
rect 254452 379652 254458 379664
rect 255038 379652 255044 379664
rect 255096 379652 255102 379704
rect 256050 379652 256056 379704
rect 256108 379692 256114 379704
rect 256510 379692 256516 379704
rect 256108 379664 256516 379692
rect 256108 379652 256114 379664
rect 256510 379652 256516 379664
rect 256568 379652 256574 379704
rect 257062 379652 257068 379704
rect 257120 379692 257126 379704
rect 257798 379692 257804 379704
rect 257120 379664 257804 379692
rect 257120 379652 257126 379664
rect 257798 379652 257804 379664
rect 257856 379652 257862 379704
rect 258046 379692 258074 379732
rect 263229 379729 263241 379732
rect 263275 379729 263287 379763
rect 263229 379723 263287 379729
rect 263428 379692 263456 379800
rect 267734 379788 267740 379800
rect 267792 379788 267798 379840
rect 263505 379763 263563 379769
rect 263505 379729 263517 379763
rect 263551 379760 263563 379763
rect 268010 379760 268016 379772
rect 263551 379732 268016 379760
rect 263551 379729 263563 379732
rect 263505 379723 263563 379729
rect 268010 379720 268016 379732
rect 268068 379720 268074 379772
rect 280522 379720 280528 379772
rect 280580 379760 280586 379772
rect 290090 379760 290096 379772
rect 280580 379732 290096 379760
rect 280580 379720 280586 379732
rect 290090 379720 290096 379732
rect 290148 379720 290154 379772
rect 258046 379664 263456 379692
rect 264422 379652 264428 379704
rect 264480 379692 264486 379704
rect 264882 379692 264888 379704
rect 264480 379664 264888 379692
rect 264480 379652 264486 379664
rect 264882 379652 264888 379664
rect 264940 379652 264946 379704
rect 265526 379652 265532 379704
rect 265584 379692 265590 379704
rect 299474 379692 299480 379704
rect 265584 379664 299480 379692
rect 265584 379652 265590 379664
rect 299474 379652 299480 379664
rect 299532 379652 299538 379704
rect 235902 379584 235908 379636
rect 235960 379624 235966 379636
rect 235960 379596 258074 379624
rect 235960 379584 235966 379596
rect 254946 379516 254952 379568
rect 255004 379556 255010 379568
rect 255222 379556 255228 379568
rect 255004 379528 255228 379556
rect 255004 379516 255010 379528
rect 255222 379516 255228 379528
rect 255280 379516 255286 379568
rect 258046 379556 258074 379596
rect 263318 379584 263324 379636
rect 263376 379624 263382 379636
rect 263502 379624 263508 379636
rect 263376 379596 263508 379624
rect 263376 379584 263382 379596
rect 263502 379584 263508 379596
rect 263560 379584 263566 379636
rect 266446 379624 266452 379636
rect 266188 379596 266452 379624
rect 266188 379556 266216 379596
rect 266446 379584 266452 379596
rect 266504 379584 266510 379636
rect 271782 379584 271788 379636
rect 271840 379624 271846 379636
rect 283282 379624 283288 379636
rect 271840 379596 283288 379624
rect 271840 379584 271846 379596
rect 283282 379584 283288 379596
rect 283340 379584 283346 379636
rect 258046 379528 266216 379556
rect 266262 379516 266268 379568
rect 266320 379556 266326 379568
rect 282914 379556 282920 379568
rect 266320 379528 282920 379556
rect 266320 379516 266326 379528
rect 282914 379516 282920 379528
rect 282972 379516 282978 379568
rect 234062 379380 234068 379432
rect 234120 379420 234126 379432
rect 283742 379420 283748 379432
rect 234120 379392 283748 379420
rect 234120 379380 234126 379392
rect 283742 379380 283748 379392
rect 283800 379380 283806 379432
rect 243354 379312 243360 379364
rect 243412 379352 243418 379364
rect 295978 379352 295984 379364
rect 243412 379324 295984 379352
rect 243412 379312 243418 379324
rect 295978 379312 295984 379324
rect 296036 379312 296042 379364
rect 232590 379244 232596 379296
rect 232648 379284 232654 379296
rect 285674 379284 285680 379296
rect 232648 379256 285680 379284
rect 232648 379244 232654 379256
rect 285674 379244 285680 379256
rect 285732 379244 285738 379296
rect 231210 379176 231216 379228
rect 231268 379216 231274 379228
rect 287146 379216 287152 379228
rect 231268 379188 287152 379216
rect 231268 379176 231274 379188
rect 287146 379176 287152 379188
rect 287204 379176 287210 379228
rect 248046 379108 248052 379160
rect 248104 379148 248110 379160
rect 302878 379148 302884 379160
rect 248104 379120 302884 379148
rect 248104 379108 248110 379120
rect 302878 379108 302884 379120
rect 302936 379108 302942 379160
rect 222930 379040 222936 379092
rect 222988 379080 222994 379092
rect 284294 379080 284300 379092
rect 222988 379052 284300 379080
rect 222988 379040 222994 379052
rect 284294 379040 284300 379052
rect 284352 379040 284358 379092
rect 242342 378972 242348 379024
rect 242400 379012 242406 379024
rect 304258 379012 304264 379024
rect 242400 378984 304264 379012
rect 242400 378972 242406 378984
rect 304258 378972 304264 378984
rect 304316 378972 304322 379024
rect 228450 378904 228456 378956
rect 228508 378944 228514 378956
rect 291654 378944 291660 378956
rect 228508 378916 291660 378944
rect 228508 378904 228514 378916
rect 291654 378904 291660 378916
rect 291712 378904 291718 378956
rect 245470 378836 245476 378888
rect 245528 378876 245534 378888
rect 307110 378876 307116 378888
rect 245528 378848 307116 378876
rect 245528 378836 245534 378848
rect 307110 378836 307116 378848
rect 307168 378836 307174 378888
rect 246022 378768 246028 378820
rect 246080 378808 246086 378820
rect 314010 378808 314016 378820
rect 246080 378780 314016 378808
rect 246080 378768 246086 378780
rect 314010 378768 314016 378780
rect 314068 378768 314074 378820
rect 249150 378700 249156 378752
rect 249208 378740 249214 378752
rect 318058 378740 318064 378752
rect 249208 378712 318064 378740
rect 249208 378700 249214 378712
rect 318058 378700 318064 378712
rect 318116 378700 318122 378752
rect 215938 378632 215944 378684
rect 215996 378672 216002 378684
rect 287422 378672 287428 378684
rect 215996 378644 287428 378672
rect 215996 378632 216002 378644
rect 287422 378632 287428 378644
rect 287480 378632 287486 378684
rect 213178 378564 213184 378616
rect 213236 378604 213242 378616
rect 292206 378604 292212 378616
rect 213236 378576 292212 378604
rect 213236 378564 213242 378576
rect 292206 378564 292212 378576
rect 292264 378564 292270 378616
rect 3602 378496 3608 378548
rect 3660 378536 3666 378548
rect 282178 378536 282184 378548
rect 3660 378508 282184 378536
rect 3660 378496 3666 378508
rect 282178 378496 282184 378508
rect 282236 378496 282242 378548
rect 248230 378428 248236 378480
rect 248288 378468 248294 378480
rect 580166 378468 580172 378480
rect 248288 378440 580172 378468
rect 248288 378428 248294 378440
rect 580166 378428 580172 378440
rect 580224 378428 580230 378480
rect 239674 378360 239680 378412
rect 239732 378400 239738 378412
rect 582653 378403 582711 378409
rect 582653 378400 582665 378403
rect 239732 378372 582665 378400
rect 239732 378360 239738 378372
rect 582653 378369 582665 378372
rect 582699 378369 582711 378403
rect 582653 378363 582711 378369
rect 240042 378292 240048 378344
rect 240100 378332 240106 378344
rect 582837 378335 582895 378341
rect 582837 378332 582849 378335
rect 240100 378304 582849 378332
rect 240100 378292 240106 378304
rect 582837 378301 582849 378304
rect 582883 378301 582895 378335
rect 582837 378295 582895 378301
rect 237190 378224 237196 378276
rect 237248 378264 237254 378276
rect 582469 378267 582527 378273
rect 582469 378264 582481 378267
rect 237248 378236 582481 378264
rect 237248 378224 237254 378236
rect 582469 378233 582481 378236
rect 582515 378233 582527 378267
rect 582469 378227 582527 378233
rect 237098 378156 237104 378208
rect 237156 378196 237162 378208
rect 582377 378199 582435 378205
rect 582377 378196 582389 378199
rect 237156 378168 582389 378196
rect 237156 378156 237162 378168
rect 582377 378165 582389 378168
rect 582423 378165 582435 378199
rect 582377 378159 582435 378165
rect 244918 377884 244924 377936
rect 244976 377924 244982 377936
rect 253201 377927 253259 377933
rect 253201 377924 253213 377927
rect 244976 377896 253213 377924
rect 244976 377884 244982 377896
rect 253201 377893 253213 377896
rect 253247 377893 253259 377927
rect 253201 377887 253259 377893
rect 246574 377816 246580 377868
rect 246632 377856 246638 377868
rect 300210 377856 300216 377868
rect 246632 377828 300216 377856
rect 246632 377816 246638 377828
rect 300210 377816 300216 377828
rect 300268 377816 300274 377868
rect 243906 377748 243912 377800
rect 243964 377788 243970 377800
rect 253109 377791 253167 377797
rect 253109 377788 253121 377791
rect 243964 377760 253121 377788
rect 243964 377748 243970 377760
rect 253109 377757 253121 377760
rect 253155 377757 253167 377791
rect 253109 377751 253167 377757
rect 253201 377791 253259 377797
rect 253201 377757 253213 377791
rect 253247 377788 253259 377791
rect 298830 377788 298836 377800
rect 253247 377760 298836 377788
rect 253247 377757 253259 377760
rect 253201 377751 253259 377757
rect 298830 377748 298836 377760
rect 298888 377748 298894 377800
rect 224218 377680 224224 377732
rect 224276 377720 224282 377732
rect 282914 377720 282920 377732
rect 224276 377692 282920 377720
rect 224276 377680 224282 377692
rect 282914 377680 282920 377692
rect 282972 377680 282978 377732
rect 246942 377612 246948 377664
rect 247000 377652 247006 377664
rect 253109 377655 253167 377661
rect 247000 377624 248414 377652
rect 247000 377612 247006 377624
rect 238570 377584 238576 377596
rect 238531 377556 238576 377584
rect 238570 377544 238576 377556
rect 238628 377544 238634 377596
rect 239214 377584 239220 377596
rect 239175 377556 239220 377584
rect 239214 377544 239220 377556
rect 239272 377544 239278 377596
rect 240778 377584 240784 377596
rect 240739 377556 240784 377584
rect 240778 377544 240784 377556
rect 240836 377544 240842 377596
rect 241606 377584 241612 377596
rect 241567 377556 241612 377584
rect 241606 377544 241612 377556
rect 241664 377544 241670 377596
rect 247586 377584 247592 377596
rect 247547 377556 247592 377584
rect 247586 377544 247592 377556
rect 247644 377544 247650 377596
rect 248386 377584 248414 377624
rect 253109 377621 253121 377655
rect 253155 377652 253167 377655
rect 305638 377652 305644 377664
rect 253155 377624 305644 377652
rect 253155 377621 253167 377624
rect 253109 377615 253167 377621
rect 305638 377612 305644 377624
rect 305696 377612 305702 377664
rect 309778 377584 309784 377596
rect 248386 377556 309784 377584
rect 309778 377544 309784 377556
rect 309836 377544 309842 377596
rect 3510 377476 3516 377528
rect 3568 377516 3574 377528
rect 271782 377516 271788 377528
rect 3568 377488 271788 377516
rect 3568 377476 3574 377488
rect 271782 377476 271788 377488
rect 271840 377476 271846 377528
rect 3418 377408 3424 377460
rect 3476 377448 3482 377460
rect 280522 377448 280528 377460
rect 3476 377420 280528 377448
rect 3476 377408 3482 377420
rect 280522 377408 280528 377420
rect 280580 377408 280586 377460
rect 284846 377448 284852 377460
rect 284807 377420 284852 377448
rect 284846 377408 284852 377420
rect 284904 377408 284910 377460
rect 220170 377340 220176 377392
rect 220228 377380 220234 377392
rect 285858 377380 285864 377392
rect 220228 377352 285864 377380
rect 220228 377340 220234 377352
rect 285858 377340 285864 377352
rect 285916 377340 285922 377392
rect 288526 377380 288532 377392
rect 288487 377352 288532 377380
rect 288526 377340 288532 377352
rect 288584 377340 288590 377392
rect 290642 377380 290648 377392
rect 290603 377352 290648 377380
rect 290642 377340 290648 377352
rect 290700 377340 290706 377392
rect 293218 377340 293224 377392
rect 293276 377340 293282 377392
rect 226978 377272 226984 377324
rect 227036 377312 227042 377324
rect 293236 377312 293264 377340
rect 227036 377284 293264 377312
rect 227036 377272 227042 377284
rect 247589 377247 247647 377253
rect 247589 377213 247601 377247
rect 247635 377244 247647 377247
rect 316678 377244 316684 377256
rect 247635 377216 316684 377244
rect 247635 377213 247647 377216
rect 247589 377207 247647 377213
rect 316678 377204 316684 377216
rect 316736 377204 316742 377256
rect 214558 377136 214564 377188
rect 214616 377176 214622 377188
rect 290645 377179 290703 377185
rect 290645 377176 290657 377179
rect 214616 377148 290657 377176
rect 214616 377136 214622 377148
rect 290645 377145 290657 377148
rect 290691 377145 290703 377179
rect 290645 377139 290703 377145
rect 209038 377068 209044 377120
rect 209096 377108 209102 377120
rect 284849 377111 284907 377117
rect 284849 377108 284861 377111
rect 209096 377080 284861 377108
rect 209096 377068 209102 377080
rect 284849 377077 284861 377080
rect 284895 377077 284907 377111
rect 284849 377071 284907 377077
rect 4798 377000 4804 377052
rect 4856 377040 4862 377052
rect 288529 377043 288587 377049
rect 288529 377040 288541 377043
rect 4856 377012 288541 377040
rect 4856 377000 4862 377012
rect 288529 377009 288541 377012
rect 288575 377009 288587 377043
rect 288529 377003 288587 377009
rect 240781 376975 240839 376981
rect 240781 376941 240793 376975
rect 240827 376972 240839 376975
rect 583021 376975 583079 376981
rect 583021 376972 583033 376975
rect 240827 376944 583033 376972
rect 240827 376941 240839 376944
rect 240781 376935 240839 376941
rect 583021 376941 583033 376944
rect 583067 376941 583079 376975
rect 583021 376935 583079 376941
rect 241609 376907 241667 376913
rect 241609 376873 241621 376907
rect 241655 376904 241667 376907
rect 583113 376907 583171 376913
rect 583113 376904 583125 376907
rect 241655 376876 583125 376904
rect 241655 376873 241667 376876
rect 241609 376867 241667 376873
rect 583113 376873 583125 376876
rect 583159 376873 583171 376907
rect 583113 376867 583171 376873
rect 239217 376839 239275 376845
rect 239217 376805 239229 376839
rect 239263 376836 239275 376839
rect 582745 376839 582803 376845
rect 582745 376836 582757 376839
rect 239263 376808 582757 376836
rect 239263 376805 239275 376808
rect 239217 376799 239275 376805
rect 582745 376805 582757 376808
rect 582791 376805 582803 376839
rect 582745 376799 582803 376805
rect 238573 376771 238631 376777
rect 238573 376737 238585 376771
rect 238619 376768 238631 376771
rect 582561 376771 582619 376777
rect 582561 376768 582573 376771
rect 238619 376740 582573 376768
rect 238619 376737 238631 376740
rect 238573 376731 238631 376737
rect 582561 376737 582573 376740
rect 582607 376737 582619 376771
rect 582561 376731 582619 376737
rect 318058 365644 318064 365696
rect 318116 365684 318122 365696
rect 580166 365684 580172 365696
rect 318116 365656 580172 365684
rect 318116 365644 318122 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 302878 353200 302884 353252
rect 302936 353240 302942 353252
rect 580166 353240 580172 353252
rect 302936 353212 580172 353240
rect 302936 353200 302942 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 3142 346332 3148 346384
rect 3200 346372 3206 346384
rect 224218 346372 224224 346384
rect 3200 346344 224224 346372
rect 3200 346332 3206 346344
rect 224218 346332 224224 346344
rect 224276 346332 224282 346384
rect 234586 338048 247770 338076
rect 125502 337628 125508 337680
rect 125560 337668 125566 337680
rect 234586 337668 234614 338048
rect 236549 338011 236607 338017
rect 236549 337977 236561 338011
rect 236595 338008 236607 338011
rect 236595 337980 246666 338008
rect 236595 337977 236607 337980
rect 236549 337971 236607 337977
rect 246638 337952 246666 337980
rect 247742 337952 247770 338048
rect 280065 338011 280123 338017
rect 280065 338008 280077 338011
rect 276354 337980 280077 338008
rect 276354 337952 276382 337980
rect 280065 337977 280077 337980
rect 280111 337977 280123 338011
rect 280065 337971 280123 337977
rect 238984 337900 238990 337952
rect 239042 337900 239048 337952
rect 239352 337940 239358 337952
rect 239324 337900 239358 337940
rect 239410 337900 239416 337952
rect 244964 337940 244970 337952
rect 244246 337912 244970 337940
rect 234798 337832 234804 337884
rect 234856 337872 234862 337884
rect 235580 337872 235586 337884
rect 234856 337844 235586 337872
rect 234856 337832 234862 337844
rect 235580 337832 235586 337844
rect 235638 337832 235644 337884
rect 238616 337832 238622 337884
rect 238674 337832 238680 337884
rect 125560 337640 234614 337668
rect 125560 337628 125566 337640
rect 237926 337628 237932 337680
rect 237984 337668 237990 337680
rect 238634 337668 238662 337832
rect 239002 337816 239030 337900
rect 239002 337776 239036 337816
rect 239030 337764 239036 337776
rect 239088 337764 239094 337816
rect 237984 337640 238662 337668
rect 237984 337628 237990 337640
rect 239214 337628 239220 337680
rect 239272 337668 239278 337680
rect 239324 337668 239352 337900
rect 242020 337832 242026 337884
rect 242078 337832 242084 337884
rect 243216 337832 243222 337884
rect 243274 337832 243280 337884
rect 243354 337832 243360 337884
rect 243412 337832 243418 337884
rect 239272 337640 239352 337668
rect 239272 337628 239278 337640
rect 241514 337628 241520 337680
rect 241572 337668 241578 337680
rect 242038 337668 242066 337832
rect 243234 337736 243262 337832
rect 242912 337708 243262 337736
rect 242912 337680 242940 337708
rect 241572 337640 242066 337668
rect 241572 337628 241578 337640
rect 242894 337628 242900 337680
rect 242952 337628 242958 337680
rect 243078 337628 243084 337680
rect 243136 337668 243142 337680
rect 243372 337668 243400 337832
rect 243136 337640 243400 337668
rect 243136 337628 243142 337640
rect 122098 337560 122104 337612
rect 122156 337600 122162 337612
rect 236549 337603 236607 337609
rect 236549 337600 236561 337603
rect 122156 337572 236561 337600
rect 122156 337560 122162 337572
rect 236549 337569 236561 337572
rect 236595 337569 236607 337603
rect 236549 337563 236607 337569
rect 97902 337492 97908 337544
rect 97960 337532 97966 337544
rect 244246 337532 244274 337912
rect 244964 337900 244970 337912
rect 245022 337900 245028 337952
rect 246068 337900 246074 337952
rect 246126 337900 246132 337952
rect 246620 337900 246626 337952
rect 246678 337900 246684 337952
rect 247264 337900 247270 337952
rect 247322 337900 247328 337952
rect 247724 337900 247730 337952
rect 247782 337900 247788 337952
rect 251128 337900 251134 337952
rect 251186 337900 251192 337952
rect 262950 337900 262956 337952
rect 263008 337900 263014 337952
rect 263824 337900 263830 337952
rect 263882 337940 263888 337952
rect 264057 337943 264115 337949
rect 264057 337940 264069 337943
rect 263882 337912 264069 337940
rect 263882 337900 263888 337912
rect 264057 337909 264069 337912
rect 264103 337909 264115 337943
rect 264057 337903 264115 337909
rect 264192 337900 264198 337952
rect 264250 337949 264256 337952
rect 264250 337943 264299 337949
rect 264250 337909 264253 337943
rect 264287 337909 264299 337943
rect 264250 337903 264299 337909
rect 264250 337900 264256 337903
rect 264560 337900 264566 337952
rect 264618 337940 264624 337952
rect 267553 337943 267611 337949
rect 267553 337940 267565 337943
rect 264618 337912 267565 337940
rect 264618 337900 264624 337912
rect 267553 337909 267565 337912
rect 267599 337909 267611 337943
rect 267553 337903 267611 337909
rect 273441 337943 273499 337949
rect 273441 337909 273453 337943
rect 273487 337940 273499 337943
rect 274404 337940 274410 337952
rect 273487 337912 274410 337940
rect 273487 337909 273499 337912
rect 273441 337903 273499 337909
rect 274404 337900 274410 337912
rect 274462 337900 274468 337952
rect 276336 337900 276342 337952
rect 276394 337900 276400 337952
rect 276704 337900 276710 337952
rect 276762 337949 276768 337952
rect 276762 337943 276811 337949
rect 276762 337909 276765 337943
rect 276799 337909 276811 337943
rect 276762 337903 276811 337909
rect 276762 337900 276768 337903
rect 277072 337900 277078 337952
rect 277130 337940 277136 337952
rect 278593 337943 278651 337949
rect 278593 337940 278605 337943
rect 277130 337912 278605 337940
rect 277130 337900 277136 337912
rect 278593 337909 278605 337912
rect 278639 337909 278651 337943
rect 278593 337903 278651 337909
rect 280433 337943 280491 337949
rect 280433 337909 280445 337943
rect 280479 337940 280491 337943
rect 281212 337940 281218 337952
rect 280479 337912 281218 337940
rect 280479 337909 280491 337912
rect 280433 337903 280491 337909
rect 281212 337900 281218 337912
rect 281270 337900 281276 337952
rect 283650 337940 283656 337952
rect 283611 337912 283656 337940
rect 283650 337900 283656 337912
rect 283708 337900 283714 337952
rect 283972 337900 283978 337952
rect 284030 337949 284036 337952
rect 284030 337943 284079 337949
rect 284030 337909 284033 337943
rect 284067 337909 284079 337943
rect 284030 337903 284079 337909
rect 284030 337900 284036 337903
rect 290596 337900 290602 337952
rect 290654 337940 290660 337952
rect 294325 337943 294383 337949
rect 294325 337940 294337 337943
rect 290654 337912 294337 337940
rect 290654 337900 290660 337912
rect 294325 337909 294337 337912
rect 294371 337909 294383 337943
rect 294325 337903 294383 337909
rect 294460 337900 294466 337952
rect 294518 337940 294524 337952
rect 294966 337940 294972 337952
rect 294518 337912 294972 337940
rect 294518 337900 294524 337912
rect 294966 337900 294972 337912
rect 295024 337900 295030 337952
rect 245056 337813 245062 337816
rect 245013 337807 245062 337813
rect 245013 337773 245025 337807
rect 245059 337773 245062 337807
rect 245013 337767 245062 337773
rect 245056 337764 245062 337767
rect 245114 337764 245120 337816
rect 246086 337736 246114 337900
rect 246160 337832 246166 337884
rect 246218 337832 246224 337884
rect 247282 337872 247310 337900
rect 247190 337844 247310 337872
rect 245764 337708 246114 337736
rect 245764 337680 245792 337708
rect 245746 337628 245752 337680
rect 245804 337628 245810 337680
rect 246022 337628 246028 337680
rect 246080 337668 246086 337680
rect 246178 337668 246206 337832
rect 247190 337680 247218 337844
rect 247310 337764 247316 337816
rect 247368 337804 247374 337816
rect 248092 337804 248098 337816
rect 247368 337776 248098 337804
rect 247368 337764 247374 337776
rect 248092 337764 248098 337776
rect 248150 337764 248156 337816
rect 250898 337764 250904 337816
rect 250956 337764 250962 337816
rect 250916 337736 250944 337764
rect 250778 337708 250944 337736
rect 250778 337680 250806 337708
rect 246080 337640 246206 337668
rect 246080 337628 246086 337640
rect 247126 337628 247132 337680
rect 247184 337640 247218 337680
rect 247184 337628 247190 337640
rect 250714 337628 250720 337680
rect 250772 337640 250806 337680
rect 250772 337628 250778 337640
rect 250898 337628 250904 337680
rect 250956 337668 250962 337680
rect 251146 337668 251174 337900
rect 251269 337875 251327 337881
rect 251269 337841 251281 337875
rect 251315 337872 251327 337875
rect 251496 337872 251502 337884
rect 251315 337844 251502 337872
rect 251315 337841 251327 337844
rect 251269 337835 251327 337841
rect 251496 337832 251502 337844
rect 251554 337832 251560 337884
rect 251772 337832 251778 337884
rect 251830 337832 251836 337884
rect 253106 337872 253112 337884
rect 253032 337844 253112 337872
rect 251790 337680 251818 337832
rect 250956 337640 251174 337668
rect 250956 337628 250962 337640
rect 251726 337628 251732 337680
rect 251784 337640 251818 337680
rect 253032 337668 253060 337844
rect 253106 337832 253112 337844
rect 253164 337832 253170 337884
rect 253612 337832 253618 337884
rect 253670 337832 253676 337884
rect 253704 337832 253710 337884
rect 253762 337832 253768 337884
rect 256004 337832 256010 337884
rect 256062 337832 256068 337884
rect 261248 337872 261254 337884
rect 260852 337844 261254 337872
rect 253106 337696 253112 337748
rect 253164 337736 253170 337748
rect 253630 337736 253658 337832
rect 253164 337708 253658 337736
rect 253164 337696 253170 337708
rect 253382 337668 253388 337680
rect 253032 337640 253388 337668
rect 251784 337628 251790 337640
rect 253382 337628 253388 337640
rect 253440 337628 253446 337680
rect 253566 337628 253572 337680
rect 253624 337668 253630 337680
rect 253722 337668 253750 337832
rect 255636 337764 255642 337816
rect 255694 337804 255700 337816
rect 255777 337807 255835 337813
rect 255777 337804 255789 337807
rect 255694 337776 255789 337804
rect 255694 337764 255700 337776
rect 255777 337773 255789 337776
rect 255823 337773 255835 337807
rect 255777 337767 255835 337773
rect 253624 337640 253750 337668
rect 253624 337628 253630 337640
rect 255682 337628 255688 337680
rect 255740 337668 255746 337680
rect 256022 337668 256050 337832
rect 260852 337816 260880 337844
rect 261248 337832 261254 337844
rect 261306 337832 261312 337884
rect 258672 337764 258678 337816
rect 258730 337764 258736 337816
rect 260834 337764 260840 337816
rect 260892 337764 260898 337816
rect 255740 337640 256050 337668
rect 255740 337628 255746 337640
rect 257430 337628 257436 337680
rect 257488 337668 257494 337680
rect 258690 337668 258718 337764
rect 257488 337640 258718 337668
rect 262968 337668 262996 337900
rect 264790 337832 264796 337884
rect 264848 337832 264854 337884
rect 269896 337832 269902 337884
rect 269954 337872 269960 337884
rect 270129 337875 270187 337881
rect 270129 337872 270141 337875
rect 269954 337844 270141 337872
rect 269954 337832 269960 337844
rect 270129 337841 270141 337844
rect 270175 337841 270187 337875
rect 270129 337835 270187 337841
rect 270632 337832 270638 337884
rect 270690 337872 270696 337884
rect 271325 337875 271383 337881
rect 271325 337872 271337 337875
rect 270690 337844 271337 337872
rect 270690 337832 270696 337844
rect 271325 337841 271337 337844
rect 271371 337841 271383 337875
rect 271325 337835 271383 337841
rect 271460 337832 271466 337884
rect 271518 337881 271524 337884
rect 271518 337875 271567 337881
rect 271518 337841 271521 337875
rect 271555 337841 271567 337875
rect 271518 337835 271567 337841
rect 271518 337832 271524 337835
rect 272564 337832 272570 337884
rect 272622 337872 272628 337884
rect 274913 337875 274971 337881
rect 274913 337872 274925 337875
rect 272622 337844 274925 337872
rect 272622 337832 272628 337844
rect 274913 337841 274925 337844
rect 274959 337841 274971 337875
rect 274913 337835 274971 337841
rect 278176 337832 278182 337884
rect 278234 337881 278240 337884
rect 278234 337875 278283 337881
rect 278234 337841 278237 337875
rect 278271 337841 278283 337875
rect 278234 337835 278283 337841
rect 278234 337832 278240 337835
rect 280016 337832 280022 337884
rect 280074 337872 280080 337884
rect 287701 337875 287759 337881
rect 287701 337872 287713 337875
rect 280074 337844 287713 337872
rect 280074 337832 280080 337844
rect 287701 337841 287713 337844
rect 287747 337841 287759 337875
rect 287701 337835 287759 337841
rect 293632 337832 293638 337884
rect 293690 337872 293696 337884
rect 294233 337875 294291 337881
rect 294233 337872 294245 337875
rect 293690 337844 294245 337872
rect 293690 337832 293696 337844
rect 294233 337841 294245 337844
rect 294279 337841 294291 337875
rect 294233 337835 294291 337841
rect 294644 337832 294650 337884
rect 294702 337872 294708 337884
rect 294874 337872 294880 337884
rect 294702 337844 294880 337872
rect 294702 337832 294708 337844
rect 294874 337832 294880 337844
rect 294932 337832 294938 337884
rect 263042 337668 263048 337680
rect 262968 337640 263048 337668
rect 257488 337628 257494 337640
rect 263042 337628 263048 337640
rect 263100 337628 263106 337680
rect 264698 337628 264704 337680
rect 264756 337668 264762 337680
rect 264808 337668 264836 337832
rect 280936 337764 280942 337816
rect 280994 337804 281000 337816
rect 281166 337804 281172 337816
rect 280994 337776 281172 337804
rect 280994 337764 281000 337776
rect 281166 337764 281172 337776
rect 281224 337764 281230 337816
rect 284340 337764 284346 337816
rect 284398 337813 284404 337816
rect 284398 337807 284447 337813
rect 284398 337773 284401 337807
rect 284435 337773 284447 337807
rect 284398 337767 284447 337773
rect 284398 337764 284404 337767
rect 285076 337764 285082 337816
rect 285134 337804 285140 337816
rect 286045 337807 286103 337813
rect 286045 337804 286057 337807
rect 285134 337776 286057 337804
rect 285134 337764 285140 337776
rect 286045 337773 286057 337776
rect 286091 337773 286103 337807
rect 286045 337767 286103 337773
rect 286180 337764 286186 337816
rect 286238 337804 286244 337816
rect 289357 337807 289415 337813
rect 289357 337804 289369 337807
rect 286238 337776 289369 337804
rect 286238 337764 286244 337776
rect 289357 337773 289369 337776
rect 289403 337773 289415 337807
rect 289357 337767 289415 337773
rect 264756 337640 264836 337668
rect 264756 337628 264762 337640
rect 270770 337628 270776 337680
rect 270828 337668 270834 337680
rect 349154 337668 349160 337680
rect 270828 337640 349160 337668
rect 270828 337628 270834 337640
rect 349154 337628 349160 337640
rect 349212 337628 349218 337680
rect 272242 337560 272248 337612
rect 272300 337600 272306 337612
rect 360838 337600 360844 337612
rect 272300 337572 360844 337600
rect 272300 337560 272306 337572
rect 360838 337560 360844 337572
rect 360896 337560 360902 337612
rect 273438 337532 273444 337544
rect 97960 337504 244274 337532
rect 273399 337504 273444 337532
rect 97960 337492 97966 337504
rect 273438 337492 273444 337504
rect 273496 337492 273502 337544
rect 274913 337535 274971 337541
rect 274913 337501 274925 337535
rect 274959 337532 274971 337535
rect 367094 337532 367100 337544
rect 274959 337504 367100 337532
rect 274959 337501 274971 337504
rect 274913 337495 274971 337501
rect 367094 337492 367100 337504
rect 367152 337492 367158 337544
rect 91002 337424 91008 337476
rect 91060 337464 91066 337476
rect 244182 337464 244188 337476
rect 91060 337436 244188 337464
rect 91060 337424 91066 337436
rect 244182 337424 244188 337436
rect 244240 337424 244246 337476
rect 272886 337424 272892 337476
rect 272944 337464 272950 337476
rect 369854 337464 369860 337476
rect 272944 337436 369860 337464
rect 272944 337424 272950 337436
rect 369854 337424 369860 337436
rect 369912 337424 369918 337476
rect 86862 337356 86868 337408
rect 86920 337396 86926 337408
rect 243814 337396 243820 337408
rect 86920 337368 243820 337396
rect 86920 337356 86926 337368
rect 243814 337356 243820 337368
rect 243872 337356 243878 337408
rect 278958 337356 278964 337408
rect 279016 337396 279022 337408
rect 425698 337396 425704 337408
rect 279016 337368 425704 337396
rect 279016 337356 279022 337368
rect 425698 337356 425704 337368
rect 425756 337356 425762 337408
rect 81342 337288 81348 337340
rect 81400 337328 81406 337340
rect 242894 337328 242900 337340
rect 81400 337300 242900 337328
rect 81400 337288 81406 337300
rect 242894 337288 242900 337300
rect 242952 337288 242958 337340
rect 279050 337288 279056 337340
rect 279108 337328 279114 337340
rect 427814 337328 427820 337340
rect 279108 337300 427820 337328
rect 279108 337288 279114 337300
rect 427814 337288 427820 337300
rect 427872 337288 427878 337340
rect 70302 337220 70308 337272
rect 70360 337260 70366 337272
rect 241514 337260 241520 337272
rect 70360 337232 241520 337260
rect 70360 337220 70366 337232
rect 241514 337220 241520 337232
rect 241572 337220 241578 337272
rect 279418 337220 279424 337272
rect 279476 337260 279482 337272
rect 432046 337260 432052 337272
rect 279476 337232 432052 337260
rect 279476 337220 279482 337232
rect 432046 337220 432052 337232
rect 432104 337220 432110 337272
rect 66162 337152 66168 337204
rect 66220 337192 66226 337204
rect 241698 337192 241704 337204
rect 66220 337164 241704 337192
rect 66220 337152 66226 337164
rect 241698 337152 241704 337164
rect 241756 337152 241762 337204
rect 280430 337192 280436 337204
rect 280391 337164 280436 337192
rect 280430 337152 280436 337164
rect 280488 337152 280494 337204
rect 287701 337195 287759 337201
rect 287701 337161 287713 337195
rect 287747 337192 287759 337195
rect 436738 337192 436744 337204
rect 287747 337164 436744 337192
rect 287747 337161 287759 337164
rect 287701 337155 287759 337161
rect 436738 337152 436744 337164
rect 436796 337152 436802 337204
rect 50338 337084 50344 337136
rect 50396 337124 50402 337136
rect 239490 337124 239496 337136
rect 50396 337096 239496 337124
rect 50396 337084 50402 337096
rect 239490 337084 239496 337096
rect 239548 337084 239554 337136
rect 283282 337084 283288 337136
rect 283340 337124 283346 337136
rect 468478 337124 468484 337136
rect 283340 337096 468484 337124
rect 283340 337084 283346 337096
rect 468478 337084 468484 337096
rect 468536 337084 468542 337136
rect 48222 337016 48228 337068
rect 48280 337056 48286 337068
rect 239858 337056 239864 337068
rect 48280 337028 239864 337056
rect 48280 337016 48286 337028
rect 239858 337016 239864 337028
rect 239916 337016 239922 337068
rect 283466 337016 283472 337068
rect 283524 337056 283530 337068
rect 470594 337056 470600 337068
rect 283524 337028 470600 337056
rect 283524 337016 283530 337028
rect 470594 337016 470600 337028
rect 470652 337016 470658 337068
rect 41322 336948 41328 337000
rect 41380 336988 41386 337000
rect 239122 336988 239128 337000
rect 41380 336960 239128 336988
rect 41380 336948 41386 336960
rect 239122 336948 239128 336960
rect 239180 336948 239186 337000
rect 283653 336991 283711 336997
rect 283653 336957 283665 336991
rect 283699 336988 283711 336991
rect 472618 336988 472624 337000
rect 283699 336960 472624 336988
rect 283699 336957 283711 336960
rect 283653 336951 283711 336957
rect 472618 336948 472624 336960
rect 472676 336948 472682 337000
rect 34422 336880 34428 336932
rect 34480 336920 34486 336932
rect 238386 336920 238392 336932
rect 34480 336892 238392 336920
rect 34480 336880 34486 336892
rect 238386 336880 238392 336892
rect 238444 336880 238450 336932
rect 292942 336880 292948 336932
rect 293000 336920 293006 336932
rect 560938 336920 560944 336932
rect 293000 336892 560944 336920
rect 293000 336880 293006 336892
rect 560938 336880 560944 336892
rect 560996 336880 561002 336932
rect 29638 336812 29644 336864
rect 29696 336852 29702 336864
rect 237650 336852 237656 336864
rect 29696 336824 237656 336852
rect 29696 336812 29702 336824
rect 237650 336812 237656 336824
rect 237708 336812 237714 336864
rect 294138 336812 294144 336864
rect 294196 336852 294202 336864
rect 574094 336852 574100 336864
rect 294196 336824 574100 336852
rect 294196 336812 294202 336824
rect 574094 336812 574100 336824
rect 574152 336812 574158 336864
rect 12342 336744 12348 336796
rect 12400 336784 12406 336796
rect 236178 336784 236184 336796
rect 12400 336756 236184 336784
rect 12400 336744 12406 336756
rect 236178 336744 236184 336756
rect 236236 336744 236242 336796
rect 263520 336756 263640 336784
rect 224218 336676 224224 336728
rect 224276 336716 224282 336728
rect 251910 336716 251916 336728
rect 224276 336688 251916 336716
rect 224276 336676 224282 336688
rect 251910 336676 251916 336688
rect 251968 336676 251974 336728
rect 252005 336719 252063 336725
rect 252005 336685 252017 336719
rect 252051 336716 252063 336719
rect 253566 336716 253572 336728
rect 252051 336688 253572 336716
rect 252051 336685 252063 336688
rect 252005 336679 252063 336685
rect 253566 336676 253572 336688
rect 253624 336676 253630 336728
rect 263410 336676 263416 336728
rect 263468 336716 263474 336728
rect 263520 336716 263548 336756
rect 263468 336688 263548 336716
rect 263612 336716 263640 336756
rect 280706 336744 280712 336796
rect 280764 336784 280770 336796
rect 280890 336784 280896 336796
rect 280764 336756 280896 336784
rect 280764 336744 280770 336756
rect 280890 336744 280896 336756
rect 280948 336744 280954 336796
rect 284846 336744 284852 336796
rect 284904 336784 284910 336796
rect 285030 336784 285036 336796
rect 284904 336756 285036 336784
rect 284904 336744 284910 336756
rect 285030 336744 285036 336756
rect 285088 336744 285094 336796
rect 294966 336744 294972 336796
rect 295024 336784 295030 336796
rect 582929 336787 582987 336793
rect 582929 336784 582941 336787
rect 295024 336756 582941 336784
rect 295024 336744 295030 336756
rect 582929 336753 582941 336756
rect 582975 336753 582987 336787
rect 582929 336747 582987 336753
rect 263612 336688 264376 336716
rect 263468 336676 263474 336688
rect 239401 336651 239459 336657
rect 239401 336617 239413 336651
rect 239447 336648 239459 336651
rect 260650 336648 260656 336660
rect 239447 336620 260656 336648
rect 239447 336617 239459 336620
rect 239401 336611 239459 336617
rect 260650 336608 260656 336620
rect 260708 336608 260714 336660
rect 262306 336608 262312 336660
rect 262364 336648 262370 336660
rect 262490 336648 262496 336660
rect 262364 336620 262496 336648
rect 262364 336608 262370 336620
rect 262490 336608 262496 336620
rect 262548 336608 262554 336660
rect 233050 336540 233056 336592
rect 233108 336580 233114 336592
rect 261018 336580 261024 336592
rect 233108 336552 261024 336580
rect 233108 336540 233114 336552
rect 261018 336540 261024 336552
rect 261076 336540 261082 336592
rect 228358 336472 228364 336524
rect 228416 336512 228422 336524
rect 258074 336512 258080 336524
rect 228416 336484 258080 336512
rect 228416 336472 228422 336484
rect 258074 336472 258080 336484
rect 258132 336472 258138 336524
rect 262490 336472 262496 336524
rect 262548 336512 262554 336524
rect 263594 336512 263600 336524
rect 262548 336484 263600 336512
rect 262548 336472 262554 336484
rect 263594 336472 263600 336484
rect 263652 336472 263658 336524
rect 222838 336404 222844 336456
rect 222896 336444 222902 336456
rect 249153 336447 249211 336453
rect 222896 336416 249104 336444
rect 222896 336404 222902 336416
rect 206278 336336 206284 336388
rect 206336 336376 206342 336388
rect 248969 336379 249027 336385
rect 248969 336376 248981 336379
rect 206336 336348 248981 336376
rect 206336 336336 206342 336348
rect 248969 336345 248981 336348
rect 249015 336345 249027 336379
rect 249076 336376 249104 336416
rect 249153 336413 249165 336447
rect 249199 336444 249211 336447
rect 252554 336444 252560 336456
rect 249199 336416 252560 336444
rect 249199 336413 249211 336416
rect 249153 336407 249211 336413
rect 252554 336404 252560 336416
rect 252612 336404 252618 336456
rect 252646 336404 252652 336456
rect 252704 336444 252710 336456
rect 256142 336444 256148 336456
rect 252704 336416 256148 336444
rect 252704 336404 252710 336416
rect 256142 336404 256148 336416
rect 256200 336404 256206 336456
rect 262214 336404 262220 336456
rect 262272 336444 262278 336456
rect 263870 336444 263876 336456
rect 262272 336416 263876 336444
rect 262272 336404 262278 336416
rect 263870 336404 263876 336416
rect 263928 336404 263934 336456
rect 256970 336376 256976 336388
rect 249076 336348 256976 336376
rect 248969 336339 249027 336345
rect 256970 336336 256976 336348
rect 257028 336336 257034 336388
rect 264348 336376 264376 336688
rect 264698 336676 264704 336728
rect 264756 336716 264762 336728
rect 292485 336719 292543 336725
rect 292485 336716 292497 336719
rect 264756 336688 292497 336716
rect 264756 336676 264762 336688
rect 292485 336685 292497 336688
rect 292531 336685 292543 336719
rect 292485 336679 292543 336685
rect 292577 336719 292635 336725
rect 292577 336685 292589 336719
rect 292623 336716 292635 336719
rect 298738 336716 298744 336728
rect 292623 336688 298744 336716
rect 292623 336685 292635 336688
rect 292577 336679 292635 336685
rect 298738 336676 298744 336688
rect 298796 336676 298802 336728
rect 272610 336608 272616 336660
rect 272668 336648 272674 336660
rect 273162 336648 273168 336660
rect 272668 336620 273168 336648
rect 272668 336608 272674 336620
rect 273162 336608 273168 336620
rect 273220 336608 273226 336660
rect 273901 336651 273959 336657
rect 273901 336617 273913 336651
rect 273947 336648 273959 336651
rect 282733 336651 282791 336657
rect 282733 336648 282745 336651
rect 273947 336620 282745 336648
rect 273947 336617 273959 336620
rect 273901 336611 273959 336617
rect 282733 336617 282745 336620
rect 282779 336617 282791 336651
rect 282733 336611 282791 336617
rect 285858 336608 285864 336660
rect 285916 336648 285922 336660
rect 320818 336648 320824 336660
rect 285916 336620 320824 336648
rect 285916 336608 285922 336620
rect 320818 336608 320824 336620
rect 320876 336608 320882 336660
rect 266538 336540 266544 336592
rect 266596 336580 266602 336592
rect 285122 336580 285128 336592
rect 266596 336552 285128 336580
rect 266596 336540 266602 336552
rect 285122 336540 285128 336552
rect 285180 336540 285186 336592
rect 286962 336540 286968 336592
rect 287020 336580 287026 336592
rect 322198 336580 322204 336592
rect 287020 336552 322204 336580
rect 287020 336540 287026 336552
rect 322198 336540 322204 336552
rect 322256 336540 322262 336592
rect 265802 336472 265808 336524
rect 265860 336512 265866 336524
rect 273901 336515 273959 336521
rect 273901 336512 273913 336515
rect 265860 336484 273913 336512
rect 265860 336472 265866 336484
rect 273901 336481 273913 336484
rect 273947 336481 273959 336515
rect 273901 336475 273959 336481
rect 273993 336515 274051 336521
rect 273993 336481 274005 336515
rect 274039 336512 274051 336515
rect 286594 336512 286600 336524
rect 274039 336484 286600 336512
rect 274039 336481 274051 336484
rect 273993 336475 274051 336481
rect 286594 336472 286600 336484
rect 286652 336472 286658 336524
rect 287330 336472 287336 336524
rect 287388 336512 287394 336524
rect 294785 336515 294843 336521
rect 294785 336512 294797 336515
rect 287388 336484 294797 336512
rect 287388 336472 287394 336484
rect 294785 336481 294797 336484
rect 294831 336481 294843 336515
rect 294785 336475 294843 336481
rect 294877 336515 294935 336521
rect 294877 336481 294889 336515
rect 294923 336512 294935 336515
rect 323670 336512 323676 336524
rect 294923 336484 323676 336512
rect 294923 336481 294935 336484
rect 294877 336475 294935 336481
rect 323670 336472 323676 336484
rect 323728 336472 323734 336524
rect 265434 336404 265440 336456
rect 265492 336444 265498 336456
rect 282457 336447 282515 336453
rect 282457 336444 282469 336447
rect 265492 336416 282469 336444
rect 265492 336404 265498 336416
rect 282457 336413 282469 336416
rect 282503 336413 282515 336447
rect 282457 336407 282515 336413
rect 282638 336404 282644 336456
rect 282696 336444 282702 336456
rect 282822 336444 282828 336456
rect 282696 336416 282828 336444
rect 282696 336404 282702 336416
rect 282822 336404 282828 336416
rect 282880 336404 282886 336456
rect 283193 336447 283251 336453
rect 283193 336413 283205 336447
rect 283239 336444 283251 336447
rect 289078 336444 289084 336456
rect 283239 336416 289084 336444
rect 283239 336413 283251 336416
rect 283193 336407 283251 336413
rect 289078 336404 289084 336416
rect 289136 336404 289142 336456
rect 289265 336447 289323 336453
rect 289265 336413 289277 336447
rect 289311 336444 289323 336447
rect 331858 336444 331864 336456
rect 289311 336416 331864 336444
rect 289311 336413 289323 336416
rect 289265 336407 289323 336413
rect 331858 336404 331864 336416
rect 331916 336404 331922 336456
rect 277486 336376 277492 336388
rect 264348 336348 277492 336376
rect 277486 336336 277492 336348
rect 277544 336336 277550 336388
rect 278041 336379 278099 336385
rect 278041 336345 278053 336379
rect 278087 336376 278099 336379
rect 323578 336376 323584 336388
rect 278087 336348 282592 336376
rect 278087 336345 278099 336348
rect 278041 336339 278099 336345
rect 204898 336268 204904 336320
rect 204956 336308 204962 336320
rect 249245 336311 249303 336317
rect 249245 336308 249257 336311
rect 204956 336280 249257 336308
rect 204956 336268 204962 336280
rect 249245 336277 249257 336280
rect 249291 336277 249303 336311
rect 249245 336271 249303 336277
rect 266906 336268 266912 336320
rect 266964 336308 266970 336320
rect 273073 336311 273131 336317
rect 273073 336308 273085 336311
rect 266964 336280 273085 336308
rect 266964 336268 266970 336280
rect 273073 336277 273085 336280
rect 273119 336277 273131 336311
rect 273073 336271 273131 336277
rect 273806 336268 273812 336320
rect 273864 336308 273870 336320
rect 274358 336308 274364 336320
rect 273864 336280 274364 336308
rect 273864 336268 273870 336280
rect 274358 336268 274364 336280
rect 274416 336268 274422 336320
rect 277394 336268 277400 336320
rect 277452 336308 277458 336320
rect 282365 336311 282423 336317
rect 282365 336308 282377 336311
rect 277452 336280 282377 336308
rect 277452 336268 277458 336280
rect 282365 336277 282377 336280
rect 282411 336277 282423 336311
rect 282564 336308 282592 336348
rect 282748 336348 323584 336376
rect 282748 336308 282776 336348
rect 323578 336336 323584 336348
rect 323636 336336 323642 336388
rect 282564 336280 282776 336308
rect 282825 336311 282883 336317
rect 282365 336271 282423 336277
rect 282825 336277 282837 336311
rect 282871 336308 282883 336311
rect 335998 336308 336004 336320
rect 282871 336280 336004 336308
rect 282871 336277 282883 336280
rect 282825 336271 282883 336277
rect 335998 336268 336004 336280
rect 336056 336268 336062 336320
rect 197998 336200 198004 336252
rect 198056 336240 198062 336252
rect 249061 336243 249119 336249
rect 249061 336240 249073 336243
rect 198056 336212 249073 336240
rect 198056 336200 198062 336212
rect 249061 336209 249073 336212
rect 249107 336209 249119 336243
rect 252005 336243 252063 336249
rect 252005 336240 252017 336243
rect 249061 336203 249119 336209
rect 249168 336212 252017 336240
rect 202138 336132 202144 336184
rect 202196 336172 202202 336184
rect 248969 336175 249027 336181
rect 248969 336172 248981 336175
rect 202196 336144 248981 336172
rect 202196 336132 202202 336144
rect 248969 336141 248981 336144
rect 249015 336141 249027 336175
rect 248969 336135 249027 336141
rect 196618 336064 196624 336116
rect 196676 336104 196682 336116
rect 249168 336104 249196 336212
rect 252005 336209 252017 336212
rect 252051 336209 252063 336243
rect 252005 336203 252063 336209
rect 252554 336200 252560 336252
rect 252612 336240 252618 336252
rect 258810 336240 258816 336252
rect 252612 336212 258816 336240
rect 252612 336200 252618 336212
rect 258810 336200 258816 336212
rect 258868 336200 258874 336252
rect 265158 336200 265164 336252
rect 265216 336240 265222 336252
rect 273165 336243 273223 336249
rect 273165 336240 273177 336243
rect 265216 336212 273177 336240
rect 265216 336200 265222 336212
rect 273165 336209 273177 336212
rect 273211 336209 273223 336243
rect 273165 336203 273223 336209
rect 280065 336243 280123 336249
rect 280065 336209 280077 336243
rect 280111 336240 280123 336243
rect 376018 336240 376024 336252
rect 280111 336212 376024 336240
rect 280111 336209 280123 336212
rect 280065 336203 280123 336209
rect 376018 336200 376024 336212
rect 376076 336200 376082 336252
rect 251266 336132 251272 336184
rect 251324 336172 251330 336184
rect 251450 336172 251456 336184
rect 251324 336144 251456 336172
rect 251324 336132 251330 336144
rect 251450 336132 251456 336144
rect 251508 336132 251514 336184
rect 251818 336132 251824 336184
rect 251876 336172 251882 336184
rect 260006 336172 260012 336184
rect 251876 336144 260012 336172
rect 251876 336132 251882 336144
rect 260006 336132 260012 336144
rect 260064 336132 260070 336184
rect 268654 336132 268660 336184
rect 268712 336172 268718 336184
rect 278041 336175 278099 336181
rect 278041 336172 278053 336175
rect 268712 336144 278053 336172
rect 268712 336132 268718 336144
rect 278041 336141 278053 336144
rect 278087 336141 278099 336175
rect 278041 336135 278099 336141
rect 278593 336175 278651 336181
rect 278593 336141 278605 336175
rect 278639 336172 278651 336175
rect 393958 336172 393964 336184
rect 278639 336144 393964 336172
rect 278639 336141 278651 336144
rect 278593 336135 278651 336141
rect 393958 336132 393964 336144
rect 394016 336132 394022 336184
rect 196676 336076 249196 336104
rect 249245 336107 249303 336113
rect 196676 336064 196682 336076
rect 249245 336073 249257 336107
rect 249291 336104 249303 336107
rect 254026 336104 254032 336116
rect 249291 336076 254032 336104
rect 249291 336073 249303 336076
rect 249245 336067 249303 336073
rect 254026 336064 254032 336076
rect 254084 336064 254090 336116
rect 263042 336064 263048 336116
rect 263100 336104 263106 336116
rect 284294 336104 284300 336116
rect 263100 336076 284300 336104
rect 263100 336064 263106 336076
rect 284294 336064 284300 336076
rect 284352 336064 284358 336116
rect 285950 336064 285956 336116
rect 286008 336104 286014 336116
rect 289265 336107 289323 336113
rect 289265 336104 289277 336107
rect 286008 336076 289277 336104
rect 286008 336064 286014 336076
rect 289265 336073 289277 336076
rect 289311 336073 289323 336107
rect 289265 336067 289323 336073
rect 289357 336107 289415 336113
rect 289357 336073 289369 336107
rect 289403 336104 289415 336107
rect 497458 336104 497464 336116
rect 289403 336076 497464 336104
rect 289403 336073 289415 336076
rect 289357 336067 289415 336073
rect 497458 336064 497464 336076
rect 497516 336064 497522 336116
rect 195238 335996 195244 336048
rect 195296 336036 195302 336048
rect 249061 336039 249119 336045
rect 249061 336036 249073 336039
rect 195296 336008 249073 336036
rect 195296 335996 195302 336008
rect 249061 336005 249073 336008
rect 249107 336005 249119 336039
rect 249061 335999 249119 336005
rect 249153 336039 249211 336045
rect 249153 336005 249165 336039
rect 249199 336036 249211 336039
rect 253014 336036 253020 336048
rect 249199 336008 253020 336036
rect 249199 336005 249211 336008
rect 249153 335999 249211 336005
rect 253014 335996 253020 336008
rect 253072 335996 253078 336048
rect 265250 335996 265256 336048
rect 265308 336036 265314 336048
rect 272886 336036 272892 336048
rect 265308 336008 272892 336036
rect 265308 335996 265314 336008
rect 272886 335996 272892 336008
rect 272944 335996 272950 336048
rect 286962 336036 286968 336048
rect 273088 336008 286968 336036
rect 231762 335928 231768 335980
rect 231820 335968 231826 335980
rect 260374 335968 260380 335980
rect 231820 335940 260380 335968
rect 231820 335928 231826 335940
rect 260374 335928 260380 335940
rect 260432 335928 260438 335980
rect 266078 335928 266084 335980
rect 266136 335968 266142 335980
rect 272797 335971 272855 335977
rect 272797 335968 272809 335971
rect 266136 335940 272809 335968
rect 266136 335928 266142 335940
rect 272797 335937 272809 335940
rect 272843 335937 272855 335971
rect 272797 335931 272855 335937
rect 231118 335860 231124 335912
rect 231176 335900 231182 335912
rect 248785 335903 248843 335909
rect 248785 335900 248797 335903
rect 231176 335872 248797 335900
rect 231176 335860 231182 335872
rect 248785 335869 248797 335872
rect 248831 335869 248843 335903
rect 248785 335863 248843 335869
rect 249061 335903 249119 335909
rect 249061 335869 249073 335903
rect 249107 335900 249119 335903
rect 254762 335900 254768 335912
rect 249107 335872 254768 335900
rect 249107 335869 249119 335872
rect 249061 335863 249119 335869
rect 254762 335860 254768 335872
rect 254820 335860 254826 335912
rect 262950 335860 262956 335912
rect 263008 335900 263014 335912
rect 266998 335900 267004 335912
rect 263008 335872 267004 335900
rect 263008 335860 263014 335872
rect 266998 335860 267004 335872
rect 267056 335860 267062 335912
rect 232498 335792 232504 335844
rect 232556 335832 232562 335844
rect 248877 335835 248935 335841
rect 248877 335832 248889 335835
rect 232556 335804 248889 335832
rect 232556 335792 232562 335804
rect 248877 335801 248889 335804
rect 248923 335801 248935 335835
rect 248877 335795 248935 335801
rect 248969 335835 249027 335841
rect 248969 335801 248981 335835
rect 249015 335832 249027 335835
rect 255130 335832 255136 335844
rect 249015 335804 255136 335832
rect 249015 335801 249027 335804
rect 248969 335795 249027 335801
rect 255130 335792 255136 335804
rect 255188 335792 255194 335844
rect 264057 335835 264115 335841
rect 264057 335801 264069 335835
rect 264103 335832 264115 335835
rect 272886 335832 272892 335844
rect 264103 335804 272892 335832
rect 264103 335801 264115 335804
rect 264057 335795 264115 335801
rect 272886 335792 272892 335804
rect 272944 335792 272950 335844
rect 233970 335724 233976 335776
rect 234028 335764 234034 335776
rect 258442 335764 258448 335776
rect 234028 335736 258448 335764
rect 234028 335724 234034 335736
rect 258442 335724 258448 335736
rect 258500 335724 258506 335776
rect 272797 335767 272855 335773
rect 272797 335733 272809 335767
rect 272843 335764 272855 335767
rect 273088 335764 273116 336008
rect 286962 335996 286968 336008
rect 287020 335996 287026 336048
rect 287698 335996 287704 336048
rect 287756 336036 287762 336048
rect 294877 336039 294935 336045
rect 294877 336036 294889 336039
rect 287756 336008 294889 336036
rect 287756 335996 287762 336008
rect 294877 336005 294889 336008
rect 294923 336005 294935 336039
rect 294877 335999 294935 336005
rect 294966 335996 294972 336048
rect 295024 336036 295030 336048
rect 295242 336036 295248 336048
rect 295024 336008 295248 336036
rect 295024 335996 295030 336008
rect 295242 335996 295248 336008
rect 295300 335996 295306 336048
rect 297361 336039 297419 336045
rect 297361 336005 297373 336039
rect 297407 336036 297419 336039
rect 522298 336036 522304 336048
rect 297407 336008 522304 336036
rect 297407 336005 297419 336008
rect 297361 335999 297419 336005
rect 522298 335996 522304 336008
rect 522356 335996 522362 336048
rect 278133 335971 278191 335977
rect 278133 335937 278145 335971
rect 278179 335968 278191 335971
rect 288529 335971 288587 335977
rect 288529 335968 288541 335971
rect 278179 335940 288541 335968
rect 278179 335937 278191 335940
rect 278133 335931 278191 335937
rect 288529 335937 288541 335940
rect 288575 335937 288587 335971
rect 288529 335931 288587 335937
rect 289538 335928 289544 335980
rect 289596 335968 289602 335980
rect 303246 335968 303252 335980
rect 289596 335940 303252 335968
rect 289596 335928 289602 335940
rect 303246 335928 303252 335940
rect 303304 335928 303310 335980
rect 273165 335903 273223 335909
rect 273165 335869 273177 335903
rect 273211 335900 273223 335903
rect 294509 335903 294567 335909
rect 294509 335900 294521 335903
rect 273211 335872 294521 335900
rect 273211 335869 273223 335872
rect 273165 335863 273223 335869
rect 294509 335869 294521 335872
rect 294555 335869 294567 335903
rect 294509 335863 294567 335869
rect 294598 335860 294604 335912
rect 294656 335900 294662 335912
rect 295150 335900 295156 335912
rect 294656 335872 295156 335900
rect 294656 335860 294662 335872
rect 295150 335860 295156 335872
rect 295208 335860 295214 335912
rect 295245 335903 295303 335909
rect 295245 335869 295257 335903
rect 295291 335900 295303 335903
rect 295702 335900 295708 335912
rect 295291 335872 295708 335900
rect 295291 335869 295303 335872
rect 295245 335863 295303 335869
rect 295702 335860 295708 335872
rect 295760 335860 295766 335912
rect 280157 335835 280215 335841
rect 280157 335801 280169 335835
rect 280203 335832 280215 335835
rect 282549 335835 282607 335841
rect 282549 335832 282561 335835
rect 280203 335804 282561 335832
rect 280203 335801 280215 335804
rect 280157 335795 280215 335801
rect 282549 335801 282561 335804
rect 282595 335801 282607 335835
rect 282549 335795 282607 335801
rect 282822 335792 282828 335844
rect 282880 335832 282886 335844
rect 287514 335832 287520 335844
rect 282880 335804 287520 335832
rect 282880 335792 282886 335804
rect 287514 335792 287520 335804
rect 287572 335792 287578 335844
rect 288066 335792 288072 335844
rect 288124 335832 288130 335844
rect 299474 335832 299480 335844
rect 288124 335804 299480 335832
rect 288124 335792 288130 335804
rect 299474 335792 299480 335804
rect 299532 335792 299538 335844
rect 304166 335832 304172 335844
rect 302206 335804 304172 335832
rect 272843 335736 273116 335764
rect 273257 335767 273315 335773
rect 272843 335733 272855 335736
rect 272797 335727 272855 335733
rect 273257 335733 273269 335767
rect 273303 335764 273315 335767
rect 276934 335764 276940 335776
rect 273303 335736 276940 335764
rect 273303 335733 273315 335736
rect 273257 335727 273315 335733
rect 276934 335724 276940 335736
rect 276992 335724 276998 335776
rect 278314 335724 278320 335776
rect 278372 335764 278378 335776
rect 283193 335767 283251 335773
rect 283193 335764 283205 335767
rect 278372 335736 283205 335764
rect 278372 335724 278378 335736
rect 283193 335733 283205 335736
rect 283239 335733 283251 335767
rect 283193 335727 283251 335733
rect 283285 335767 283343 335773
rect 283285 335733 283297 335767
rect 283331 335764 283343 335767
rect 285214 335764 285220 335776
rect 283331 335736 285220 335764
rect 283331 335733 283343 335736
rect 283285 335727 283343 335733
rect 285214 335724 285220 335736
rect 285272 335724 285278 335776
rect 285490 335764 285496 335776
rect 285451 335736 285496 335764
rect 285490 335724 285496 335736
rect 285548 335724 285554 335776
rect 286502 335724 286508 335776
rect 286560 335764 286566 335776
rect 296622 335764 296628 335776
rect 286560 335736 296628 335764
rect 286560 335724 286566 335736
rect 296622 335724 296628 335736
rect 296680 335724 296686 335776
rect 233878 335656 233884 335708
rect 233936 335696 233942 335708
rect 249153 335699 249211 335705
rect 233936 335668 249104 335696
rect 233936 335656 233942 335668
rect 234430 335588 234436 335640
rect 234488 335628 234494 335640
rect 248969 335631 249027 335637
rect 248969 335628 248981 335631
rect 234488 335600 248981 335628
rect 234488 335588 234494 335600
rect 248969 335597 248981 335600
rect 249015 335597 249027 335631
rect 249076 335628 249104 335668
rect 249153 335665 249165 335699
rect 249199 335696 249211 335699
rect 259178 335696 259184 335708
rect 249199 335668 259184 335696
rect 249199 335665 249211 335668
rect 249153 335659 249211 335665
rect 259178 335656 259184 335668
rect 259236 335656 259242 335708
rect 269574 335656 269580 335708
rect 269632 335696 269638 335708
rect 272981 335699 273039 335705
rect 272981 335696 272993 335699
rect 269632 335668 272993 335696
rect 269632 335656 269638 335668
rect 272981 335665 272993 335668
rect 273027 335665 273039 335699
rect 272981 335659 273039 335665
rect 273073 335699 273131 335705
rect 273073 335665 273085 335699
rect 273119 335696 273131 335699
rect 273993 335699 274051 335705
rect 273993 335696 274005 335699
rect 273119 335668 274005 335696
rect 273119 335665 273131 335668
rect 273073 335659 273131 335665
rect 273993 335665 274005 335668
rect 274039 335665 274051 335699
rect 273993 335659 274051 335665
rect 278194 335668 278452 335696
rect 254394 335628 254400 335640
rect 249076 335600 254400 335628
rect 248969 335591 249027 335597
rect 254394 335588 254400 335600
rect 254452 335588 254458 335640
rect 266722 335588 266728 335640
rect 266780 335628 266786 335640
rect 278194 335628 278222 335668
rect 266780 335600 278222 335628
rect 278424 335628 278452 335668
rect 278498 335656 278504 335708
rect 278556 335696 278562 335708
rect 278682 335696 278688 335708
rect 278556 335668 278688 335696
rect 278556 335656 278562 335668
rect 278682 335656 278688 335668
rect 278740 335656 278746 335708
rect 279510 335656 279516 335708
rect 279568 335696 279574 335708
rect 279694 335696 279700 335708
rect 279568 335668 279700 335696
rect 279568 335656 279574 335668
rect 279694 335656 279700 335668
rect 279752 335656 279758 335708
rect 281353 335699 281411 335705
rect 281353 335665 281365 335699
rect 281399 335696 281411 335699
rect 283101 335699 283159 335705
rect 281399 335668 282684 335696
rect 281399 335665 281411 335668
rect 281353 335659 281411 335665
rect 278424 335600 282592 335628
rect 266780 335588 266786 335600
rect 230474 335520 230480 335572
rect 230532 335560 230538 335572
rect 252278 335560 252284 335572
rect 230532 335532 252284 335560
rect 230532 335520 230538 335532
rect 252278 335520 252284 335532
rect 252336 335520 252342 335572
rect 253842 335520 253848 335572
rect 253900 335560 253906 335572
rect 262306 335560 262312 335572
rect 253900 335532 262312 335560
rect 253900 335520 253906 335532
rect 262306 335520 262312 335532
rect 262364 335520 262370 335572
rect 268010 335520 268016 335572
rect 268068 335560 268074 335572
rect 278133 335563 278191 335569
rect 278133 335560 278145 335563
rect 268068 335532 278145 335560
rect 268068 335520 268074 335532
rect 278133 335529 278145 335532
rect 278179 335529 278191 335563
rect 278133 335523 278191 335529
rect 278314 335520 278320 335572
rect 278372 335560 278378 335572
rect 278372 335532 281580 335560
rect 278372 335520 278378 335532
rect 233142 335452 233148 335504
rect 233200 335492 233206 335504
rect 248877 335495 248935 335501
rect 233200 335464 247908 335492
rect 233200 335452 233206 335464
rect 233418 335384 233424 335436
rect 233476 335424 233482 335436
rect 247880 335424 247908 335464
rect 248877 335461 248889 335495
rect 248923 335492 248935 335495
rect 257338 335492 257344 335504
rect 248923 335464 257344 335492
rect 248923 335461 248935 335464
rect 248877 335455 248935 335461
rect 257338 335452 257344 335464
rect 257396 335452 257402 335504
rect 260098 335452 260104 335504
rect 260156 335492 260162 335504
rect 261294 335492 261300 335504
rect 260156 335464 261300 335492
rect 260156 335452 260162 335464
rect 261294 335452 261300 335464
rect 261352 335452 261358 335504
rect 262766 335452 262772 335504
rect 262824 335492 262830 335504
rect 263502 335492 263508 335504
rect 262824 335464 263508 335492
rect 262824 335452 262830 335464
rect 263502 335452 263508 335464
rect 263560 335452 263566 335504
rect 269758 335452 269764 335504
rect 269816 335492 269822 335504
rect 270126 335492 270132 335504
rect 269816 335464 270132 335492
rect 269816 335452 269822 335464
rect 270126 335452 270132 335464
rect 270184 335452 270190 335504
rect 271966 335452 271972 335504
rect 272024 335492 272030 335504
rect 272886 335492 272892 335504
rect 272024 335464 272892 335492
rect 272024 335452 272030 335464
rect 272886 335452 272892 335464
rect 272944 335452 272950 335504
rect 272981 335495 273039 335501
rect 272981 335461 272993 335495
rect 273027 335492 273039 335495
rect 273257 335495 273315 335501
rect 273257 335492 273269 335495
rect 273027 335464 273269 335492
rect 273027 335461 273039 335464
rect 272981 335455 273039 335461
rect 273257 335461 273269 335464
rect 273303 335461 273315 335495
rect 273257 335455 273315 335461
rect 273346 335452 273352 335504
rect 273404 335492 273410 335504
rect 273404 335464 274588 335492
rect 273404 335452 273410 335464
rect 251269 335427 251327 335433
rect 251269 335424 251281 335427
rect 233476 335396 244274 335424
rect 247880 335396 251281 335424
rect 233476 335384 233482 335396
rect 231670 335316 231676 335368
rect 231728 335356 231734 335368
rect 239401 335359 239459 335365
rect 239401 335356 239413 335359
rect 231728 335328 239413 335356
rect 231728 335316 231734 335328
rect 239401 335325 239413 335328
rect 239447 335325 239459 335359
rect 244246 335356 244274 335396
rect 251269 335393 251281 335396
rect 251315 335393 251327 335427
rect 251269 335387 251327 335393
rect 251361 335427 251419 335433
rect 251361 335393 251373 335427
rect 251407 335424 251419 335427
rect 253290 335424 253296 335436
rect 251407 335396 253296 335424
rect 251407 335393 251419 335396
rect 251361 335387 251419 335393
rect 253290 335384 253296 335396
rect 253348 335384 253354 335436
rect 257706 335424 257712 335436
rect 253906 335396 257712 335424
rect 248693 335359 248751 335365
rect 248693 335356 248705 335359
rect 244246 335328 248705 335356
rect 239401 335319 239459 335325
rect 248693 335325 248705 335328
rect 248739 335325 248751 335359
rect 248693 335319 248751 335325
rect 248785 335359 248843 335365
rect 248785 335325 248797 335359
rect 248831 335356 248843 335359
rect 253906 335356 253934 335396
rect 257706 335384 257712 335396
rect 257764 335384 257770 335436
rect 260650 335384 260656 335436
rect 260708 335424 260714 335436
rect 261754 335424 261760 335436
rect 260708 335396 261760 335424
rect 260708 335384 260714 335396
rect 261754 335384 261760 335396
rect 261812 335384 261818 335436
rect 262582 335384 262588 335436
rect 262640 335424 262646 335436
rect 263410 335424 263416 335436
rect 262640 335396 263416 335424
rect 262640 335384 262646 335396
rect 263410 335384 263416 335396
rect 263468 335384 263474 335436
rect 265066 335384 265072 335436
rect 265124 335424 265130 335436
rect 265802 335424 265808 335436
rect 265124 335396 265808 335424
rect 265124 335384 265130 335396
rect 265802 335384 265808 335396
rect 265860 335384 265866 335436
rect 268654 335384 268660 335436
rect 268712 335424 268718 335436
rect 269022 335424 269028 335436
rect 268712 335396 269028 335424
rect 268712 335384 268718 335396
rect 269022 335384 269028 335396
rect 269080 335384 269086 335436
rect 271322 335384 271328 335436
rect 271380 335424 271386 335436
rect 271690 335424 271696 335436
rect 271380 335396 271696 335424
rect 271380 335384 271386 335396
rect 271690 335384 271696 335396
rect 271748 335384 271754 335436
rect 272334 335384 272340 335436
rect 272392 335424 272398 335436
rect 273070 335424 273076 335436
rect 272392 335396 273076 335424
rect 272392 335384 272398 335396
rect 273070 335384 273076 335396
rect 273128 335384 273134 335436
rect 248831 335328 253934 335356
rect 248831 335325 248843 335328
rect 248785 335319 248843 335325
rect 254854 335316 254860 335368
rect 254912 335356 254918 335368
rect 255774 335356 255780 335368
rect 254912 335328 255780 335356
rect 254912 335316 254918 335328
rect 255774 335316 255780 335328
rect 255832 335316 255838 335368
rect 258718 335316 258724 335368
rect 258776 335356 258782 335368
rect 259730 335356 259736 335368
rect 258776 335328 259736 335356
rect 258776 335316 258782 335328
rect 259730 335316 259736 335328
rect 259788 335316 259794 335368
rect 261110 335316 261116 335368
rect 261168 335356 261174 335368
rect 261846 335356 261852 335368
rect 261168 335328 261852 335356
rect 261168 335316 261174 335328
rect 261846 335316 261852 335328
rect 261904 335316 261910 335368
rect 266630 335316 266636 335368
rect 266688 335356 266694 335368
rect 267090 335356 267096 335368
rect 266688 335328 267096 335356
rect 266688 335316 266694 335328
rect 267090 335316 267096 335328
rect 267148 335316 267154 335368
rect 267274 335316 267280 335368
rect 267332 335356 267338 335368
rect 267826 335356 267832 335368
rect 267332 335328 267832 335356
rect 267332 335316 267338 335328
rect 267826 335316 267832 335328
rect 267884 335316 267890 335368
rect 268194 335316 268200 335368
rect 268252 335356 268258 335368
rect 268252 335328 268700 335356
rect 268252 335316 268258 335328
rect 151722 335248 151728 335300
rect 151780 335288 151786 335300
rect 250438 335288 250444 335300
rect 151780 335260 250444 335288
rect 151780 335248 151786 335260
rect 250438 335248 250444 335260
rect 250496 335248 250502 335300
rect 147582 335180 147588 335232
rect 147640 335220 147646 335232
rect 250070 335220 250076 335232
rect 147640 335192 250076 335220
rect 147640 335180 147646 335192
rect 250070 335180 250076 335192
rect 250128 335180 250134 335232
rect 262122 335180 262128 335232
rect 262180 335220 262186 335232
rect 262858 335220 262864 335232
rect 262180 335192 262864 335220
rect 262180 335180 262186 335192
rect 262858 335180 262864 335192
rect 262916 335180 262922 335232
rect 268672 335220 268700 335328
rect 268746 335316 268752 335368
rect 268804 335356 268810 335368
rect 268930 335356 268936 335368
rect 268804 335328 268936 335356
rect 268804 335316 268810 335328
rect 268930 335316 268936 335328
rect 268988 335316 268994 335368
rect 270494 335316 270500 335368
rect 270552 335356 270558 335368
rect 270954 335356 270960 335368
rect 270552 335328 270960 335356
rect 270552 335316 270558 335328
rect 270954 335316 270960 335328
rect 271012 335316 271018 335368
rect 271230 335316 271236 335368
rect 271288 335356 271294 335368
rect 271506 335356 271512 335368
rect 271288 335328 271512 335356
rect 271288 335316 271294 335328
rect 271506 335316 271512 335328
rect 271564 335316 271570 335368
rect 271874 335356 271880 335368
rect 271708 335328 271880 335356
rect 271708 335300 271736 335328
rect 271874 335316 271880 335328
rect 271932 335316 271938 335368
rect 273622 335316 273628 335368
rect 273680 335356 273686 335368
rect 274082 335356 274088 335368
rect 273680 335328 274088 335356
rect 273680 335316 273686 335328
rect 274082 335316 274088 335328
rect 274140 335316 274146 335368
rect 274560 335356 274588 335464
rect 277670 335452 277676 335504
rect 277728 335492 277734 335504
rect 278498 335492 278504 335504
rect 277728 335464 278504 335492
rect 277728 335452 277734 335464
rect 278498 335452 278504 335464
rect 278556 335452 278562 335504
rect 280157 335495 280215 335501
rect 280157 335492 280169 335495
rect 279068 335464 280169 335492
rect 275186 335384 275192 335436
rect 275244 335424 275250 335436
rect 275244 335396 276520 335424
rect 275244 335384 275250 335396
rect 274468 335328 274588 335356
rect 274468 335300 274496 335328
rect 274634 335316 274640 335368
rect 274692 335356 274698 335368
rect 275462 335356 275468 335368
rect 274692 335328 275468 335356
rect 274692 335316 274698 335328
rect 275462 335316 275468 335328
rect 275520 335316 275526 335368
rect 275922 335316 275928 335368
rect 275980 335356 275986 335368
rect 275980 335328 276428 335356
rect 275980 335316 275986 335328
rect 271690 335248 271696 335300
rect 271748 335248 271754 335300
rect 274450 335248 274456 335300
rect 274508 335248 274514 335300
rect 268746 335220 268752 335232
rect 268672 335192 268752 335220
rect 268746 335180 268752 335192
rect 268804 335180 268810 335232
rect 276400 335220 276428 335328
rect 276492 335288 276520 335396
rect 276750 335384 276756 335436
rect 276808 335424 276814 335436
rect 277302 335424 277308 335436
rect 276808 335396 277308 335424
rect 276808 335384 276814 335396
rect 277302 335384 277308 335396
rect 277360 335384 277366 335436
rect 279068 335424 279096 335464
rect 280157 335461 280169 335464
rect 280203 335461 280215 335495
rect 280157 335455 280215 335461
rect 278516 335396 279096 335424
rect 276952 335328 278084 335356
rect 276952 335288 276980 335328
rect 276492 335260 276980 335288
rect 278056 335288 278084 335328
rect 278130 335316 278136 335368
rect 278188 335356 278194 335368
rect 278406 335356 278412 335368
rect 278188 335328 278412 335356
rect 278188 335316 278194 335328
rect 278406 335316 278412 335328
rect 278464 335316 278470 335368
rect 278516 335288 278544 335396
rect 279142 335384 279148 335436
rect 279200 335424 279206 335436
rect 279878 335424 279884 335436
rect 279200 335396 279884 335424
rect 279200 335384 279206 335396
rect 279878 335384 279884 335396
rect 279936 335384 279942 335436
rect 280798 335384 280804 335436
rect 280856 335424 280862 335436
rect 281442 335424 281448 335436
rect 280856 335396 281448 335424
rect 280856 335384 280862 335396
rect 281442 335384 281448 335396
rect 281500 335384 281506 335436
rect 278774 335316 278780 335368
rect 278832 335356 278838 335368
rect 279510 335356 279516 335368
rect 278832 335328 279516 335356
rect 278832 335316 278838 335328
rect 279510 335316 279516 335328
rect 279568 335316 279574 335368
rect 281552 335356 281580 335532
rect 281552 335328 282132 335356
rect 278056 335260 278544 335288
rect 282104 335288 282132 335328
rect 282178 335316 282184 335368
rect 282236 335356 282242 335368
rect 282454 335356 282460 335368
rect 282236 335328 282460 335356
rect 282236 335316 282242 335328
rect 282454 335316 282460 335328
rect 282512 335316 282518 335368
rect 282564 335356 282592 335600
rect 282656 335560 282684 335668
rect 283101 335665 283113 335699
rect 283147 335696 283159 335699
rect 286321 335699 286379 335705
rect 286321 335696 286333 335699
rect 283147 335668 286333 335696
rect 283147 335665 283159 335668
rect 283101 335659 283159 335665
rect 286321 335665 286333 335668
rect 286367 335665 286379 335699
rect 286321 335659 286379 335665
rect 288802 335656 288808 335708
rect 288860 335696 288866 335708
rect 292393 335699 292451 335705
rect 292393 335696 292405 335699
rect 288860 335668 292405 335696
rect 288860 335656 288866 335668
rect 292393 335665 292405 335668
rect 292439 335665 292451 335699
rect 292393 335659 292451 335665
rect 292758 335656 292764 335708
rect 292816 335696 292822 335708
rect 302206 335696 302234 335804
rect 304166 335792 304172 335804
rect 304224 335792 304230 335844
rect 292816 335668 302234 335696
rect 292816 335656 292822 335668
rect 282822 335588 282828 335640
rect 282880 335628 282886 335640
rect 282880 335600 288434 335628
rect 282880 335588 282886 335600
rect 283285 335563 283343 335569
rect 283285 335560 283297 335563
rect 282656 335532 283297 335560
rect 283285 335529 283297 335532
rect 283331 335529 283343 335563
rect 285490 335560 285496 335572
rect 283285 335523 283343 335529
rect 283392 335532 285496 335560
rect 282641 335495 282699 335501
rect 282641 335461 282653 335495
rect 282687 335492 282699 335495
rect 283392 335492 283420 335532
rect 285490 335520 285496 335532
rect 285548 335520 285554 335572
rect 287238 335520 287244 335572
rect 287296 335560 287302 335572
rect 287974 335560 287980 335572
rect 287296 335532 287980 335560
rect 287296 335520 287302 335532
rect 287974 335520 287980 335532
rect 288032 335520 288038 335572
rect 284386 335492 284392 335504
rect 282687 335464 283420 335492
rect 283484 335464 284392 335492
rect 282687 335461 282699 335464
rect 282641 335455 282699 335461
rect 282733 335427 282791 335433
rect 282733 335393 282745 335427
rect 282779 335424 282791 335427
rect 283484 335424 283512 335464
rect 284386 335452 284392 335464
rect 284444 335452 284450 335504
rect 284478 335452 284484 335504
rect 284536 335492 284542 335504
rect 285398 335492 285404 335504
rect 284536 335464 285404 335492
rect 284536 335452 284542 335464
rect 285398 335452 285404 335464
rect 285456 335452 285462 335504
rect 287606 335452 287612 335504
rect 287664 335492 287670 335504
rect 288066 335492 288072 335504
rect 287664 335464 288072 335492
rect 287664 335452 287670 335464
rect 288066 335452 288072 335464
rect 288124 335452 288130 335504
rect 285674 335424 285680 335436
rect 282779 335396 283512 335424
rect 284128 335396 285680 335424
rect 282779 335393 282791 335396
rect 282733 335387 282791 335393
rect 283101 335359 283159 335365
rect 283101 335356 283113 335359
rect 282564 335328 283113 335356
rect 283101 335325 283113 335328
rect 283147 335325 283159 335359
rect 284128 335356 284156 335396
rect 285674 335384 285680 335396
rect 285732 335384 285738 335436
rect 286318 335424 286324 335436
rect 286279 335396 286324 335424
rect 286318 335384 286324 335396
rect 286376 335384 286382 335436
rect 287238 335384 287244 335436
rect 287296 335424 287302 335436
rect 287882 335424 287888 335436
rect 287296 335396 287888 335424
rect 287296 335384 287302 335396
rect 287882 335384 287888 335396
rect 287940 335384 287946 335436
rect 283101 335319 283159 335325
rect 283852 335328 284156 335356
rect 282104 335260 282914 335288
rect 281353 335223 281411 335229
rect 281353 335220 281365 335223
rect 276400 335192 281365 335220
rect 281353 335189 281365 335192
rect 281399 335189 281411 335223
rect 282886 335220 282914 335260
rect 283852 335220 283880 335328
rect 284662 335316 284668 335368
rect 284720 335356 284726 335368
rect 285398 335356 285404 335368
rect 284720 335328 285404 335356
rect 284720 335316 284726 335328
rect 285398 335316 285404 335328
rect 285456 335316 285462 335368
rect 285766 335316 285772 335368
rect 285824 335356 285830 335368
rect 286870 335356 286876 335368
rect 285824 335328 286876 335356
rect 285824 335316 285830 335328
rect 286870 335316 286876 335328
rect 286928 335316 286934 335368
rect 287698 335316 287704 335368
rect 287756 335356 287762 335368
rect 288250 335356 288256 335368
rect 287756 335328 288256 335356
rect 287756 335316 287762 335328
rect 288250 335316 288256 335328
rect 288308 335316 288314 335368
rect 288406 335288 288434 335600
rect 289170 335588 289176 335640
rect 289228 335628 289234 335640
rect 294049 335631 294107 335637
rect 294049 335628 294061 335631
rect 289228 335600 294061 335628
rect 289228 335588 289234 335600
rect 294049 335597 294061 335600
rect 294095 335597 294107 335631
rect 294049 335591 294107 335597
rect 294141 335631 294199 335637
rect 294141 335597 294153 335631
rect 294187 335628 294199 335631
rect 296530 335628 296536 335640
rect 294187 335600 296536 335628
rect 294187 335597 294199 335600
rect 294141 335591 294199 335597
rect 296530 335588 296536 335600
rect 296588 335588 296594 335640
rect 288529 335563 288587 335569
rect 288529 335529 288541 335563
rect 288575 335560 288587 335563
rect 292577 335563 292635 335569
rect 292577 335560 292589 335563
rect 288575 335532 292589 335560
rect 288575 335529 288587 335532
rect 288529 335523 288587 335529
rect 292577 335529 292589 335532
rect 292623 335529 292635 335563
rect 292577 335523 292635 335529
rect 292669 335563 292727 335569
rect 292669 335529 292681 335563
rect 292715 335560 292727 335563
rect 294785 335563 294843 335569
rect 294785 335560 294797 335563
rect 292715 335532 294797 335560
rect 292715 335529 292727 335532
rect 292669 335523 292727 335529
rect 294785 335529 294797 335532
rect 294831 335529 294843 335563
rect 294785 335523 294843 335529
rect 294874 335520 294880 335572
rect 294932 335560 294938 335572
rect 295242 335560 295248 335572
rect 294932 335532 295248 335560
rect 294932 335520 294938 335532
rect 295242 335520 295248 335532
rect 295300 335520 295306 335572
rect 295337 335563 295395 335569
rect 295337 335529 295349 335563
rect 295383 335560 295395 335563
rect 298186 335560 298192 335572
rect 295383 335532 298192 335560
rect 295383 335529 295395 335532
rect 295337 335523 295395 335529
rect 298186 335520 298192 335532
rect 298244 335520 298250 335572
rect 288618 335452 288624 335504
rect 288676 335492 288682 335504
rect 289446 335492 289452 335504
rect 288676 335464 289452 335492
rect 288676 335452 288682 335464
rect 289446 335452 289452 335464
rect 289504 335452 289510 335504
rect 289906 335452 289912 335504
rect 289964 335492 289970 335504
rect 292393 335495 292451 335501
rect 289964 335464 292298 335492
rect 289964 335452 289970 335464
rect 288986 335384 288992 335436
rect 289044 335424 289050 335436
rect 289538 335424 289544 335436
rect 289044 335396 289544 335424
rect 289044 335384 289050 335396
rect 289538 335384 289544 335396
rect 289596 335384 289602 335436
rect 292270 335424 292298 335464
rect 292393 335461 292405 335495
rect 292439 335492 292451 335495
rect 297361 335495 297419 335501
rect 297361 335492 297373 335495
rect 292439 335464 297373 335492
rect 292439 335461 292451 335464
rect 292393 335455 292451 335461
rect 297361 335461 297373 335464
rect 297407 335461 297419 335495
rect 297361 335455 297419 335461
rect 294141 335427 294199 335433
rect 294141 335424 294153 335427
rect 292270 335396 294153 335424
rect 294141 335393 294153 335396
rect 294187 335393 294199 335427
rect 294141 335387 294199 335393
rect 294230 335384 294236 335436
rect 294288 335424 294294 335436
rect 294874 335424 294880 335436
rect 294288 335396 294880 335424
rect 294288 335384 294294 335396
rect 294874 335384 294880 335396
rect 294932 335384 294938 335436
rect 294969 335427 295027 335433
rect 294969 335393 294981 335427
rect 295015 335424 295027 335427
rect 295426 335424 295432 335436
rect 295015 335396 295432 335424
rect 295015 335393 295027 335396
rect 294969 335387 295027 335393
rect 295426 335384 295432 335396
rect 295484 335384 295490 335436
rect 288894 335316 288900 335368
rect 288952 335356 288958 335368
rect 289354 335356 289360 335368
rect 288952 335328 289360 335356
rect 288952 335316 288958 335328
rect 289354 335316 289360 335328
rect 289412 335316 289418 335368
rect 290090 335316 290096 335368
rect 290148 335356 290154 335368
rect 290918 335356 290924 335368
rect 290148 335328 290924 335356
rect 290148 335316 290154 335328
rect 290918 335316 290924 335328
rect 290976 335316 290982 335368
rect 291746 335316 291752 335368
rect 291804 335356 291810 335368
rect 292114 335356 292120 335368
rect 291804 335328 292120 335356
rect 291804 335316 291810 335328
rect 292114 335316 292120 335328
rect 292172 335316 292178 335368
rect 292209 335359 292267 335365
rect 292209 335325 292221 335359
rect 292255 335356 292267 335359
rect 292574 335356 292580 335368
rect 292255 335328 292580 335356
rect 292255 335325 292267 335328
rect 292209 335319 292267 335325
rect 292574 335316 292580 335328
rect 292632 335316 292638 335368
rect 292666 335316 292672 335368
rect 292724 335356 292730 335368
rect 293862 335356 293868 335368
rect 292724 335328 293868 335356
rect 292724 335316 292730 335328
rect 293862 335316 293868 335328
rect 293920 335316 293926 335368
rect 294049 335359 294107 335365
rect 294049 335325 294061 335359
rect 294095 335356 294107 335359
rect 294693 335359 294751 335365
rect 294693 335356 294705 335359
rect 294095 335328 294705 335356
rect 294095 335325 294107 335328
rect 294049 335319 294107 335325
rect 294693 335325 294705 335328
rect 294739 335325 294751 335359
rect 294693 335319 294751 335325
rect 294782 335316 294788 335368
rect 294840 335356 294846 335368
rect 295150 335356 295156 335368
rect 294840 335328 295156 335356
rect 294840 335316 294846 335328
rect 295150 335316 295156 335328
rect 295208 335316 295214 335368
rect 295245 335359 295303 335365
rect 295245 335325 295257 335359
rect 295291 335356 295303 335359
rect 296346 335356 296352 335368
rect 295291 335328 296352 335356
rect 295291 335325 295303 335328
rect 295245 335319 295303 335325
rect 296346 335316 296352 335328
rect 296404 335316 296410 335368
rect 295061 335291 295119 335297
rect 288406 335260 294644 335288
rect 282886 335192 283880 335220
rect 285493 335223 285551 335229
rect 281353 335183 281411 335189
rect 285493 335189 285505 335223
rect 285539 335220 285551 335223
rect 292209 335223 292267 335229
rect 292209 335220 292221 335223
rect 285539 335192 292221 335220
rect 285539 335189 285551 335192
rect 285493 335183 285551 335189
rect 292209 335189 292221 335192
rect 292255 335189 292267 335223
rect 292209 335183 292267 335189
rect 292485 335223 292543 335229
rect 292485 335189 292497 335223
rect 292531 335220 292543 335223
rect 292669 335223 292727 335229
rect 292669 335220 292681 335223
rect 292531 335192 292681 335220
rect 292531 335189 292543 335192
rect 292485 335183 292543 335189
rect 292669 335189 292681 335192
rect 292715 335189 292727 335223
rect 294616 335220 294644 335260
rect 295061 335257 295073 335291
rect 295107 335288 295119 335291
rect 387794 335288 387800 335300
rect 295107 335260 387800 335288
rect 295107 335257 295119 335260
rect 295061 335251 295119 335257
rect 387794 335248 387800 335260
rect 387852 335248 387858 335300
rect 394694 335220 394700 335232
rect 294616 335192 394700 335220
rect 292669 335183 292727 335189
rect 394694 335180 394700 335192
rect 394752 335180 394758 335232
rect 144822 335112 144828 335164
rect 144880 335152 144886 335164
rect 249702 335152 249708 335164
rect 144880 335124 249708 335152
rect 144880 335112 144886 335124
rect 249702 335112 249708 335124
rect 249760 335112 249766 335164
rect 277762 335112 277768 335164
rect 277820 335152 277826 335164
rect 414658 335152 414664 335164
rect 277820 335124 414664 335152
rect 277820 335112 277826 335124
rect 414658 335112 414664 335124
rect 414716 335112 414722 335164
rect 126882 335044 126888 335096
rect 126940 335084 126946 335096
rect 234522 335084 234528 335096
rect 126940 335056 234528 335084
rect 126940 335044 126946 335056
rect 234522 335044 234528 335056
rect 234580 335044 234586 335096
rect 249334 335084 249340 335096
rect 244246 335056 249340 335084
rect 140682 334976 140688 335028
rect 140740 335016 140746 335028
rect 244246 335016 244274 335056
rect 249334 335044 249340 335056
rect 249392 335044 249398 335096
rect 279602 335044 279608 335096
rect 279660 335084 279666 335096
rect 432598 335084 432604 335096
rect 279660 335056 432604 335084
rect 279660 335044 279666 335056
rect 432598 335044 432604 335056
rect 432656 335044 432662 335096
rect 140740 334988 244274 335016
rect 248693 335019 248751 335025
rect 140740 334976 140746 334988
rect 248693 334985 248705 335019
rect 248739 335016 248751 335019
rect 251361 335019 251419 335025
rect 251361 335016 251373 335019
rect 248739 334988 251373 335016
rect 248739 334985 248751 334988
rect 248693 334979 248751 334985
rect 251361 334985 251373 334988
rect 251407 334985 251419 335019
rect 251361 334979 251419 334985
rect 263962 334976 263968 335028
rect 264020 335016 264026 335028
rect 264790 335016 264796 335028
rect 264020 334988 264796 335016
rect 264020 334976 264026 334988
rect 264790 334976 264796 334988
rect 264848 334976 264854 335028
rect 284754 334976 284760 335028
rect 284812 335016 284818 335028
rect 290001 335019 290059 335025
rect 284812 334988 289906 335016
rect 284812 334976 284818 334988
rect 137278 334908 137284 334960
rect 137336 334948 137342 334960
rect 248966 334948 248972 334960
rect 137336 334920 248972 334948
rect 137336 334908 137342 334920
rect 248966 334908 248972 334920
rect 249024 334908 249030 334960
rect 289878 334948 289906 334988
rect 290001 334985 290013 335019
rect 290047 335016 290059 335019
rect 480254 335016 480260 335028
rect 290047 334988 480260 335016
rect 290047 334985 290059 334988
rect 290001 334979 290059 334985
rect 480254 334976 480260 334988
rect 480312 334976 480318 335028
rect 483014 334948 483020 334960
rect 289878 334920 483020 334948
rect 483014 334908 483020 334920
rect 483072 334908 483078 334960
rect 133782 334840 133788 334892
rect 133840 334880 133846 334892
rect 248598 334880 248604 334892
rect 133840 334852 248604 334880
rect 133840 334840 133846 334852
rect 248598 334840 248604 334852
rect 248656 334840 248662 334892
rect 286045 334883 286103 334889
rect 286045 334849 286057 334883
rect 286091 334880 286103 334883
rect 487154 334880 487160 334892
rect 286091 334852 487160 334880
rect 286091 334849 286103 334852
rect 286045 334843 286103 334849
rect 487154 334840 487160 334852
rect 487212 334840 487218 334892
rect 128998 334772 129004 334824
rect 129056 334812 129062 334824
rect 247954 334812 247960 334824
rect 129056 334784 247960 334812
rect 129056 334772 129062 334784
rect 247954 334772 247960 334784
rect 248012 334772 248018 334824
rect 287514 334772 287520 334824
rect 287572 334812 287578 334824
rect 295061 334815 295119 334821
rect 295061 334812 295073 334815
rect 287572 334784 295073 334812
rect 287572 334772 287578 334784
rect 295061 334781 295073 334784
rect 295107 334781 295119 334815
rect 295061 334775 295119 334781
rect 296622 334772 296628 334824
rect 296680 334812 296686 334824
rect 500954 334812 500960 334824
rect 296680 334784 500960 334812
rect 296680 334772 296686 334784
rect 500954 334772 500960 334784
rect 501012 334772 501018 334824
rect 87598 334704 87604 334756
rect 87656 334744 87662 334756
rect 243630 334744 243636 334756
rect 87656 334716 243636 334744
rect 87656 334704 87662 334716
rect 243630 334704 243636 334716
rect 243688 334704 243694 334756
rect 257338 334704 257344 334756
rect 257396 334744 257402 334756
rect 260006 334744 260012 334756
rect 257396 334716 260012 334744
rect 257396 334704 257402 334716
rect 260006 334704 260012 334716
rect 260064 334704 260070 334756
rect 282086 334704 282092 334756
rect 282144 334744 282150 334756
rect 282362 334744 282368 334756
rect 282144 334716 282368 334744
rect 282144 334704 282150 334716
rect 282362 334704 282368 334716
rect 282420 334704 282426 334756
rect 284386 334704 284392 334756
rect 284444 334744 284450 334756
rect 299382 334744 299388 334756
rect 284444 334716 299388 334744
rect 284444 334704 284450 334716
rect 299382 334704 299388 334716
rect 299440 334704 299446 334756
rect 299474 334704 299480 334756
rect 299532 334744 299538 334756
rect 514754 334744 514760 334756
rect 299532 334716 514760 334744
rect 299532 334704 299538 334716
rect 514754 334704 514760 334716
rect 514812 334704 514818 334756
rect 52362 334636 52368 334688
rect 52420 334676 52426 334688
rect 240226 334676 240232 334688
rect 52420 334648 240232 334676
rect 52420 334636 52426 334648
rect 240226 334636 240232 334648
rect 240284 334636 240290 334688
rect 273254 334636 273260 334688
rect 273312 334676 273318 334688
rect 273312 334648 282914 334676
rect 273312 334636 273318 334648
rect 17862 334568 17868 334620
rect 17920 334608 17926 334620
rect 236638 334608 236644 334620
rect 17920 334580 236644 334608
rect 17920 334568 17926 334580
rect 236638 334568 236644 334580
rect 236696 334568 236702 334620
rect 237466 334568 237472 334620
rect 237524 334608 237530 334620
rect 237742 334608 237748 334620
rect 237524 334580 237748 334608
rect 237524 334568 237530 334580
rect 237742 334568 237748 334580
rect 237800 334568 237806 334620
rect 239122 334568 239128 334620
rect 239180 334608 239186 334620
rect 239674 334608 239680 334620
rect 239180 334580 239680 334608
rect 239180 334568 239186 334580
rect 239674 334568 239680 334580
rect 239732 334568 239738 334620
rect 242986 334568 242992 334620
rect 243044 334608 243050 334620
rect 243446 334608 243452 334620
rect 243044 334580 243452 334608
rect 243044 334568 243050 334580
rect 243446 334568 243452 334580
rect 243504 334568 243510 334620
rect 244918 334568 244924 334620
rect 244976 334608 244982 334620
rect 245194 334608 245200 334620
rect 244976 334580 245200 334608
rect 244976 334568 244982 334580
rect 245194 334568 245200 334580
rect 245252 334568 245258 334620
rect 246390 334568 246396 334620
rect 246448 334608 246454 334620
rect 246574 334608 246580 334620
rect 246448 334580 246580 334608
rect 246448 334568 246454 334580
rect 246574 334568 246580 334580
rect 246632 334568 246638 334620
rect 251634 334568 251640 334620
rect 251692 334608 251698 334620
rect 252462 334608 252468 334620
rect 251692 334580 252468 334608
rect 251692 334568 251698 334580
rect 252462 334568 252468 334580
rect 252520 334568 252526 334620
rect 252830 334568 252836 334620
rect 252888 334608 252894 334620
rect 253750 334608 253756 334620
rect 252888 334580 253756 334608
rect 252888 334568 252894 334580
rect 253750 334568 253756 334580
rect 253808 334568 253814 334620
rect 258350 334568 258356 334620
rect 258408 334608 258414 334620
rect 259362 334608 259368 334620
rect 258408 334580 259368 334608
rect 258408 334568 258414 334580
rect 259362 334568 259368 334580
rect 259420 334568 259426 334620
rect 260006 334568 260012 334620
rect 260064 334608 260070 334620
rect 260742 334608 260748 334620
rect 260064 334580 260748 334608
rect 260064 334568 260070 334580
rect 260742 334568 260748 334580
rect 260800 334568 260806 334620
rect 273622 334568 273628 334620
rect 273680 334608 273686 334620
rect 273990 334608 273996 334620
rect 273680 334580 273996 334608
rect 273680 334568 273686 334580
rect 273990 334568 273996 334580
rect 274048 334568 274054 334620
rect 282086 334568 282092 334620
rect 282144 334608 282150 334620
rect 282730 334608 282736 334620
rect 282144 334580 282736 334608
rect 282144 334568 282150 334580
rect 282730 334568 282736 334580
rect 282788 334568 282794 334620
rect 155218 334500 155224 334552
rect 155276 334540 155282 334552
rect 250806 334540 250812 334552
rect 155276 334512 250812 334540
rect 155276 334500 155282 334512
rect 250806 334500 250812 334512
rect 250864 334500 250870 334552
rect 271322 334540 271328 334552
rect 271283 334512 271328 334540
rect 271322 334500 271328 334512
rect 271380 334500 271386 334552
rect 275554 334500 275560 334552
rect 275612 334540 275618 334552
rect 275830 334540 275836 334552
rect 275612 334512 275836 334540
rect 275612 334500 275618 334512
rect 275830 334500 275836 334512
rect 275888 334500 275894 334552
rect 282886 334540 282914 334648
rect 285490 334636 285496 334688
rect 285548 334676 285554 334688
rect 295334 334676 295340 334688
rect 285548 334648 295340 334676
rect 285548 334636 285554 334648
rect 295334 334636 295340 334648
rect 295392 334636 295398 334688
rect 296530 334636 296536 334688
rect 296588 334676 296594 334688
rect 532694 334676 532700 334688
rect 296588 334648 532700 334676
rect 296588 334636 296594 334648
rect 532694 334636 532700 334648
rect 532752 334636 532758 334688
rect 284389 334611 284447 334617
rect 284389 334577 284401 334611
rect 284435 334608 284447 334611
rect 289909 334611 289967 334617
rect 289909 334608 289921 334611
rect 284435 334580 289921 334608
rect 284435 334577 284447 334580
rect 284389 334571 284447 334577
rect 289909 334577 289921 334580
rect 289955 334577 289967 334611
rect 289909 334571 289967 334577
rect 289998 334568 290004 334620
rect 290056 334608 290062 334620
rect 535454 334608 535460 334620
rect 290056 334580 535460 334608
rect 290056 334568 290062 334580
rect 535454 334568 535460 334580
rect 535512 334568 535518 334620
rect 371878 334540 371884 334552
rect 282886 334512 371884 334540
rect 371878 334500 371884 334512
rect 371936 334500 371942 334552
rect 158622 334432 158628 334484
rect 158680 334472 158686 334484
rect 250898 334472 250904 334484
rect 158680 334444 250904 334472
rect 158680 334432 158686 334444
rect 250898 334432 250904 334444
rect 250956 334432 250962 334484
rect 271046 334432 271052 334484
rect 271104 334472 271110 334484
rect 351914 334472 351920 334484
rect 271104 334444 351920 334472
rect 271104 334432 271110 334444
rect 351914 334432 351920 334444
rect 351972 334432 351978 334484
rect 161382 334364 161388 334416
rect 161440 334404 161446 334416
rect 233142 334404 233148 334416
rect 161440 334376 233148 334404
rect 161440 334364 161446 334376
rect 233142 334364 233148 334376
rect 233200 334364 233206 334416
rect 252554 334404 252560 334416
rect 234586 334376 252560 334404
rect 169662 334296 169668 334348
rect 169720 334336 169726 334348
rect 230474 334336 230480 334348
rect 169720 334308 230480 334336
rect 169720 334296 169726 334308
rect 230474 334296 230480 334308
rect 230532 334296 230538 334348
rect 233234 334296 233240 334348
rect 233292 334336 233298 334348
rect 234586 334336 234614 334376
rect 252554 334364 252560 334376
rect 252612 334364 252618 334416
rect 262398 334364 262404 334416
rect 262456 334404 262462 334416
rect 263410 334404 263416 334416
rect 262456 334376 263416 334404
rect 262456 334364 262462 334376
rect 263410 334364 263416 334376
rect 263468 334364 263474 334416
rect 263778 334364 263784 334416
rect 263836 334404 263842 334416
rect 264238 334404 264244 334416
rect 263836 334376 264244 334404
rect 263836 334364 263842 334376
rect 264238 334364 264244 334376
rect 264296 334364 264302 334416
rect 269206 334364 269212 334416
rect 269264 334404 269270 334416
rect 333974 334404 333980 334416
rect 269264 334376 333980 334404
rect 269264 334364 269270 334376
rect 333974 334364 333980 334376
rect 334032 334364 334038 334416
rect 233292 334308 234614 334336
rect 233292 334296 233298 334308
rect 268378 334296 268384 334348
rect 268436 334336 268442 334348
rect 324314 334336 324320 334348
rect 268436 334308 324320 334336
rect 268436 334296 268442 334308
rect 324314 334296 324320 334308
rect 324372 334296 324378 334348
rect 194410 334228 194416 334280
rect 194468 334268 194474 334280
rect 254762 334268 254768 334280
rect 194468 334240 254768 334268
rect 194468 334228 194474 334240
rect 254762 334228 254768 334240
rect 254820 334228 254826 334280
rect 267550 334228 267556 334280
rect 267608 334268 267614 334280
rect 316034 334268 316040 334280
rect 267608 334240 316040 334268
rect 267608 334228 267614 334240
rect 316034 334228 316040 334240
rect 316092 334228 316098 334280
rect 212442 334160 212448 334212
rect 212500 334200 212506 334212
rect 256786 334200 256792 334212
rect 212500 334172 256792 334200
rect 212500 334160 212506 334172
rect 256786 334160 256792 334172
rect 256844 334160 256850 334212
rect 267182 334160 267188 334212
rect 267240 334200 267246 334212
rect 313274 334200 313280 334212
rect 267240 334172 313280 334200
rect 267240 334160 267246 334172
rect 313274 334160 313280 334172
rect 313332 334160 313338 334212
rect 220078 334092 220084 334144
rect 220136 334132 220142 334144
rect 257522 334132 257528 334144
rect 220136 334104 257528 334132
rect 220136 334092 220142 334104
rect 257522 334092 257528 334104
rect 257580 334092 257586 334144
rect 286594 334092 286600 334144
rect 286652 334132 286658 334144
rect 309134 334132 309140 334144
rect 286652 334104 309140 334132
rect 286652 334092 286658 334104
rect 309134 334092 309140 334104
rect 309192 334092 309198 334144
rect 227622 334024 227628 334076
rect 227680 334064 227686 334076
rect 258258 334064 258264 334076
rect 227680 334036 258264 334064
rect 227680 334024 227686 334036
rect 258258 334024 258264 334036
rect 258316 334024 258322 334076
rect 285122 334024 285128 334076
rect 285180 334064 285186 334076
rect 306374 334064 306380 334076
rect 285180 334036 306380 334064
rect 285180 334024 285186 334036
rect 306374 334024 306380 334036
rect 306432 334024 306438 334076
rect 230382 333956 230388 334008
rect 230440 333996 230446 334008
rect 258534 333996 258540 334008
rect 230440 333968 258540 333996
rect 230440 333956 230446 333968
rect 258534 333956 258540 333968
rect 258592 333956 258598 334008
rect 286962 333956 286968 334008
rect 287020 333996 287026 334008
rect 302234 333996 302240 334008
rect 287020 333968 302240 333996
rect 287020 333956 287026 333968
rect 302234 333956 302240 333968
rect 302292 333956 302298 334008
rect 187602 333888 187608 333940
rect 187660 333928 187666 333940
rect 254210 333928 254216 333940
rect 187660 333900 254216 333928
rect 187660 333888 187666 333900
rect 254210 333888 254216 333900
rect 254268 333888 254274 333940
rect 278225 333931 278283 333937
rect 278225 333897 278237 333931
rect 278271 333928 278283 333931
rect 418798 333928 418804 333940
rect 278271 333900 418804 333928
rect 278271 333897 278283 333900
rect 278225 333891 278283 333897
rect 418798 333888 418804 333900
rect 418856 333888 418862 333940
rect 166902 333820 166908 333872
rect 166960 333860 166966 333872
rect 252002 333860 252008 333872
rect 166960 333832 252008 333860
rect 166960 333820 166966 333832
rect 252002 333820 252008 333832
rect 252060 333820 252066 333872
rect 278682 333820 278688 333872
rect 278740 333860 278746 333872
rect 423674 333860 423680 333872
rect 278740 333832 423680 333860
rect 278740 333820 278746 333832
rect 423674 333820 423680 333832
rect 423732 333820 423738 333872
rect 162762 333752 162768 333804
rect 162820 333792 162826 333804
rect 251910 333792 251916 333804
rect 162820 333764 251916 333792
rect 162820 333752 162826 333764
rect 251910 333752 251916 333764
rect 251968 333752 251974 333804
rect 287330 333752 287336 333804
rect 287388 333792 287394 333804
rect 465166 333792 465172 333804
rect 287388 333764 465172 333792
rect 287388 333752 287394 333764
rect 465166 333752 465172 333764
rect 465224 333752 465230 333804
rect 144730 333684 144736 333736
rect 144788 333724 144794 333736
rect 249794 333724 249800 333736
rect 144788 333696 249800 333724
rect 144788 333684 144794 333696
rect 249794 333684 249800 333696
rect 249852 333684 249858 333736
rect 292114 333684 292120 333736
rect 292172 333724 292178 333736
rect 292482 333724 292488 333736
rect 292172 333696 292488 333724
rect 292172 333684 292178 333696
rect 292482 333684 292488 333696
rect 292540 333684 292546 333736
rect 292574 333684 292580 333736
rect 292632 333724 292638 333736
rect 489914 333724 489920 333736
rect 292632 333696 489920 333724
rect 292632 333684 292638 333696
rect 489914 333684 489920 333696
rect 489972 333684 489978 333736
rect 135162 333616 135168 333668
rect 135220 333656 135226 333668
rect 248690 333656 248696 333668
rect 135220 333628 248696 333656
rect 135220 333616 135226 333628
rect 248690 333616 248696 333628
rect 248748 333616 248754 333668
rect 265618 333616 265624 333668
rect 265676 333656 265682 333668
rect 298094 333656 298100 333668
rect 265676 333628 298100 333656
rect 265676 333616 265682 333628
rect 298094 333616 298100 333628
rect 298152 333616 298158 333668
rect 298186 333616 298192 333668
rect 298244 333656 298250 333668
rect 507854 333656 507860 333668
rect 298244 333628 507860 333656
rect 298244 333616 298250 333628
rect 507854 333616 507860 333628
rect 507912 333616 507918 333668
rect 88978 333548 88984 333600
rect 89036 333588 89042 333600
rect 243998 333588 244004 333600
rect 89036 333560 244004 333588
rect 89036 333548 89042 333560
rect 243998 333548 244004 333560
rect 244056 333548 244062 333600
rect 287054 333548 287060 333600
rect 287112 333588 287118 333600
rect 506474 333588 506480 333600
rect 287112 333560 506480 333588
rect 287112 333548 287118 333560
rect 506474 333548 506480 333560
rect 506532 333548 506538 333600
rect 83458 333480 83464 333532
rect 83516 333520 83522 333532
rect 239306 333520 239312 333532
rect 83516 333492 239312 333520
rect 83516 333480 83522 333492
rect 239306 333480 239312 333492
rect 239364 333480 239370 333532
rect 265986 333480 265992 333532
rect 266044 333520 266050 333532
rect 300118 333520 300124 333532
rect 266044 333492 300124 333520
rect 266044 333480 266050 333492
rect 300118 333480 300124 333492
rect 300176 333480 300182 333532
rect 303246 333480 303252 333532
rect 303304 333520 303310 333532
rect 529934 333520 529940 333532
rect 303304 333492 529940 333520
rect 303304 333480 303310 333492
rect 529934 333480 529940 333492
rect 529992 333480 529998 333532
rect 73062 333412 73068 333464
rect 73120 333452 73126 333464
rect 242434 333452 242440 333464
rect 73120 333424 242440 333452
rect 73120 333412 73126 333424
rect 242434 333412 242440 333424
rect 242492 333412 242498 333464
rect 288802 333412 288808 333464
rect 288860 333452 288866 333464
rect 524506 333452 524512 333464
rect 288860 333424 524512 333452
rect 288860 333412 288866 333424
rect 524506 333412 524512 333424
rect 524564 333412 524570 333464
rect 59262 333344 59268 333396
rect 59320 333384 59326 333396
rect 240962 333384 240968 333396
rect 59320 333356 240968 333384
rect 59320 333344 59326 333356
rect 240962 333344 240968 333356
rect 241020 333344 241026 333396
rect 290734 333344 290740 333396
rect 290792 333384 290798 333396
rect 542446 333384 542452 333396
rect 290792 333356 542452 333384
rect 290792 333344 290798 333356
rect 542446 333344 542452 333356
rect 542504 333344 542510 333396
rect 55122 333276 55128 333328
rect 55180 333316 55186 333328
rect 240594 333316 240600 333328
rect 55180 333288 240600 333316
rect 55180 333276 55186 333288
rect 240594 333276 240600 333288
rect 240652 333276 240658 333328
rect 280614 333276 280620 333328
rect 280672 333316 280678 333328
rect 281258 333316 281264 333328
rect 280672 333288 281264 333316
rect 280672 333276 280678 333288
rect 281258 333276 281264 333288
rect 281316 333276 281322 333328
rect 283190 333276 283196 333328
rect 283248 333316 283254 333328
rect 283742 333316 283748 333328
rect 283248 333288 283748 333316
rect 283248 333276 283254 333288
rect 283742 333276 283748 333288
rect 283800 333276 283806 333328
rect 291194 333276 291200 333328
rect 291252 333316 291258 333328
rect 292298 333316 292304 333328
rect 291252 333288 292304 333316
rect 291252 333276 291258 333288
rect 292298 333276 292304 333288
rect 292356 333276 292362 333328
rect 296438 333276 296444 333328
rect 296496 333316 296502 333328
rect 547874 333316 547880 333328
rect 296496 333288 547880 333316
rect 296496 333276 296502 333288
rect 547874 333276 547880 333288
rect 547932 333276 547938 333328
rect 22002 333208 22008 333260
rect 22060 333248 22066 333260
rect 237190 333248 237196 333260
rect 22060 333220 237196 333248
rect 22060 333208 22066 333220
rect 237190 333208 237196 333220
rect 237248 333208 237254 333260
rect 258810 333208 258816 333260
rect 258868 333248 258874 333260
rect 259822 333248 259828 333260
rect 258868 333220 259828 333248
rect 258868 333208 258874 333220
rect 259822 333208 259828 333220
rect 259880 333208 259886 333260
rect 264054 333208 264060 333260
rect 264112 333248 264118 333260
rect 264514 333248 264520 333260
rect 264112 333220 264520 333248
rect 264112 333208 264118 333220
rect 264514 333208 264520 333220
rect 264572 333208 264578 333260
rect 265526 333208 265532 333260
rect 265584 333248 265590 333260
rect 266078 333248 266084 333260
rect 265584 333220 266084 333248
rect 265584 333208 265590 333220
rect 266078 333208 266084 333220
rect 266136 333208 266142 333260
rect 272702 333208 272708 333260
rect 272760 333248 272766 333260
rect 273162 333248 273168 333260
rect 272760 333220 273168 333248
rect 272760 333208 272766 333220
rect 273162 333208 273168 333220
rect 273220 333208 273226 333260
rect 273898 333208 273904 333260
rect 273956 333248 273962 333260
rect 274174 333248 274180 333260
rect 273956 333220 274180 333248
rect 273956 333208 273962 333220
rect 274174 333208 274180 333220
rect 274232 333208 274238 333260
rect 276474 333208 276480 333260
rect 276532 333248 276538 333260
rect 277118 333248 277124 333260
rect 276532 333220 277124 333248
rect 276532 333208 276538 333220
rect 277118 333208 277124 333220
rect 277176 333208 277182 333260
rect 277578 333208 277584 333260
rect 277636 333248 277642 333260
rect 278314 333248 278320 333260
rect 277636 333220 278320 333248
rect 277636 333208 277642 333220
rect 278314 333208 278320 333220
rect 278372 333208 278378 333260
rect 280246 333208 280252 333260
rect 280304 333248 280310 333260
rect 281442 333248 281448 333260
rect 280304 333220 281448 333248
rect 280304 333208 280310 333220
rect 281442 333208 281448 333220
rect 281500 333208 281506 333260
rect 283558 333208 283564 333260
rect 283616 333248 283622 333260
rect 284018 333248 284024 333260
rect 283616 333220 284024 333248
rect 283616 333208 283622 333220
rect 284018 333208 284024 333220
rect 284076 333208 284082 333260
rect 298002 333208 298008 333260
rect 298060 333248 298066 333260
rect 568574 333248 568580 333260
rect 298060 333220 568580 333248
rect 298060 333208 298066 333220
rect 568574 333208 568580 333220
rect 568632 333208 568638 333260
rect 169570 333140 169576 333192
rect 169628 333180 169634 333192
rect 252370 333180 252376 333192
rect 169628 333152 252376 333180
rect 169628 333140 169634 333152
rect 252370 333140 252376 333152
rect 252428 333140 252434 333192
rect 276753 333183 276811 333189
rect 276753 333149 276765 333183
rect 276799 333180 276811 333183
rect 405734 333180 405740 333192
rect 276799 333152 405740 333180
rect 276799 333149 276811 333152
rect 276753 333143 276811 333149
rect 405734 333140 405740 333152
rect 405792 333140 405798 333192
rect 191742 333072 191748 333124
rect 191800 333112 191806 333124
rect 254578 333112 254584 333124
rect 191800 333084 254584 333112
rect 191800 333072 191806 333084
rect 254578 333072 254584 333084
rect 254636 333072 254642 333124
rect 282365 333115 282423 333121
rect 282365 333081 282377 333115
rect 282411 333112 282423 333115
rect 412634 333112 412640 333124
rect 282411 333084 412640 333112
rect 282411 333081 282423 333084
rect 282365 333075 282423 333081
rect 412634 333072 412640 333084
rect 412692 333072 412698 333124
rect 198642 333004 198648 333056
rect 198700 333044 198706 333056
rect 255222 333044 255228 333056
rect 198700 333016 255228 333044
rect 198700 333004 198706 333016
rect 255222 333004 255228 333016
rect 255280 333004 255286 333056
rect 285214 333004 285220 333056
rect 285272 333044 285278 333056
rect 398834 333044 398840 333056
rect 285272 333016 398840 333044
rect 285272 333004 285278 333016
rect 398834 333004 398840 333016
rect 398892 333004 398898 333056
rect 179322 332936 179328 332988
rect 179380 332976 179386 332988
rect 233418 332976 233424 332988
rect 179380 332948 233424 332976
rect 179380 332936 179386 332948
rect 233418 332936 233424 332948
rect 233476 332936 233482 332988
rect 254578 332936 254584 332988
rect 254636 332976 254642 332988
rect 259086 332976 259092 332988
rect 254636 332948 259092 332976
rect 254636 332936 254642 332948
rect 259086 332936 259092 332948
rect 259144 332936 259150 332988
rect 271509 332979 271567 332985
rect 271509 332945 271521 332979
rect 271555 332976 271567 332979
rect 353938 332976 353944 332988
rect 271555 332948 353944 332976
rect 271555 332945 271567 332948
rect 271509 332939 271567 332945
rect 353938 332936 353944 332948
rect 353996 332936 354002 332988
rect 206922 332868 206928 332920
rect 206980 332908 206986 332920
rect 252646 332908 252652 332920
rect 206980 332880 252652 332908
rect 206980 332868 206986 332880
rect 252646 332868 252652 332880
rect 252704 332868 252710 332920
rect 269298 332868 269304 332920
rect 269356 332908 269362 332920
rect 331950 332908 331956 332920
rect 269356 332880 331956 332908
rect 269356 332868 269362 332880
rect 331950 332868 331956 332880
rect 332008 332868 332014 332920
rect 210970 332800 210976 332852
rect 211028 332840 211034 332852
rect 256510 332840 256516 332852
rect 211028 332812 256516 332840
rect 211028 332800 211034 332812
rect 256510 332800 256516 332812
rect 256568 332800 256574 332852
rect 268102 332800 268108 332852
rect 268160 332840 268166 332852
rect 321554 332840 321560 332852
rect 268160 332812 321560 332840
rect 268160 332800 268166 332812
rect 321554 332800 321560 332812
rect 321612 332800 321618 332852
rect 216582 332732 216588 332784
rect 216640 332772 216646 332784
rect 257154 332772 257160 332784
rect 216640 332744 257160 332772
rect 216640 332732 216646 332744
rect 257154 332732 257160 332744
rect 257212 332732 257218 332784
rect 266906 332732 266912 332784
rect 266964 332772 266970 332784
rect 310514 332772 310520 332784
rect 266964 332744 310520 332772
rect 266964 332732 266970 332744
rect 310514 332732 310520 332744
rect 310572 332732 310578 332784
rect 223482 332664 223488 332716
rect 223540 332704 223546 332716
rect 257798 332704 257804 332716
rect 223540 332676 257804 332704
rect 223540 332664 223546 332676
rect 257798 332664 257804 332676
rect 257856 332664 257862 332716
rect 266722 332664 266728 332716
rect 266780 332704 266786 332716
rect 307018 332704 307024 332716
rect 266780 332676 307024 332704
rect 266780 332664 266786 332676
rect 307018 332664 307024 332676
rect 307076 332664 307082 332716
rect 227530 332596 227536 332648
rect 227588 332636 227594 332648
rect 258166 332636 258172 332648
rect 227588 332608 258172 332636
rect 227588 332596 227594 332608
rect 258166 332596 258172 332608
rect 258224 332596 258230 332648
rect 153102 332528 153108 332580
rect 153160 332568 153166 332580
rect 250530 332568 250536 332580
rect 153160 332540 250536 332568
rect 153160 332528 153166 332540
rect 250530 332528 250536 332540
rect 250588 332528 250594 332580
rect 284846 332528 284852 332580
rect 284904 332568 284910 332580
rect 430574 332568 430580 332580
rect 284904 332540 430580 332568
rect 284904 332528 284910 332540
rect 430574 332528 430580 332540
rect 430632 332528 430638 332580
rect 148962 332460 148968 332512
rect 149020 332500 149026 332512
rect 250162 332500 250168 332512
rect 149020 332472 250168 332500
rect 149020 332460 149026 332472
rect 250162 332460 250168 332472
rect 250220 332460 250226 332512
rect 284021 332503 284079 332509
rect 284021 332469 284033 332503
rect 284067 332500 284079 332503
rect 476114 332500 476120 332512
rect 284067 332472 476120 332500
rect 284067 332469 284079 332472
rect 284021 332463 284079 332469
rect 476114 332460 476120 332472
rect 476172 332460 476178 332512
rect 142062 332392 142068 332444
rect 142120 332432 142126 332444
rect 249426 332432 249432 332444
rect 142120 332404 249432 332432
rect 142120 332392 142126 332404
rect 249426 332392 249432 332404
rect 249484 332392 249490 332444
rect 284570 332392 284576 332444
rect 284628 332432 284634 332444
rect 481634 332432 481640 332444
rect 284628 332404 481640 332432
rect 284628 332392 284634 332404
rect 481634 332392 481640 332404
rect 481692 332392 481698 332444
rect 137922 332324 137928 332376
rect 137980 332364 137986 332376
rect 249058 332364 249064 332376
rect 137980 332336 249064 332364
rect 137980 332324 137986 332336
rect 249058 332324 249064 332336
rect 249116 332324 249122 332376
rect 285030 332324 285036 332376
rect 285088 332364 285094 332376
rect 484394 332364 484400 332376
rect 285088 332336 484400 332364
rect 285088 332324 285094 332336
rect 484394 332324 484400 332336
rect 484452 332324 484458 332376
rect 124122 332256 124128 332308
rect 124180 332296 124186 332308
rect 247586 332296 247592 332308
rect 124180 332268 247592 332296
rect 124180 332256 124186 332268
rect 247586 332256 247592 332268
rect 247644 332256 247650 332308
rect 286226 332256 286232 332308
rect 286284 332296 286290 332308
rect 499666 332296 499672 332308
rect 286284 332268 499672 332296
rect 286284 332256 286290 332268
rect 499666 332256 499672 332268
rect 499724 332256 499730 332308
rect 104802 332188 104808 332240
rect 104860 332228 104866 332240
rect 245654 332228 245660 332240
rect 104860 332200 245660 332228
rect 104860 332188 104866 332200
rect 245654 332188 245660 332200
rect 245712 332188 245718 332240
rect 287422 332188 287428 332240
rect 287480 332228 287486 332240
rect 510706 332228 510712 332240
rect 287480 332200 510712 332228
rect 287480 332188 287486 332200
rect 510706 332188 510712 332200
rect 510764 332188 510770 332240
rect 95142 332120 95148 332172
rect 95200 332160 95206 332172
rect 244642 332160 244648 332172
rect 95200 332132 244648 332160
rect 95200 332120 95206 332132
rect 244642 332120 244648 332132
rect 244700 332120 244706 332172
rect 296346 332120 296352 332172
rect 296404 332160 296410 332172
rect 525794 332160 525800 332172
rect 296404 332132 525800 332160
rect 296404 332120 296410 332132
rect 525794 332120 525800 332132
rect 525852 332120 525858 332172
rect 77202 332052 77208 332104
rect 77260 332092 77266 332104
rect 235997 332095 236055 332101
rect 235997 332092 236009 332095
rect 77260 332064 236009 332092
rect 77260 332052 77266 332064
rect 235997 332061 236009 332064
rect 236043 332061 236055 332095
rect 241330 332092 241336 332104
rect 235997 332055 236055 332061
rect 236104 332064 241336 332092
rect 62022 331984 62028 332036
rect 62080 332024 62086 332036
rect 236104 332024 236132 332064
rect 241330 332052 241336 332064
rect 241388 332052 241394 332104
rect 288526 332052 288532 332104
rect 288584 332092 288590 332104
rect 520274 332092 520280 332104
rect 288584 332064 520280 332092
rect 288584 332052 288590 332064
rect 520274 332052 520280 332064
rect 520332 332052 520338 332104
rect 239950 332024 239956 332036
rect 62080 331996 236132 332024
rect 236242 331996 239956 332024
rect 62080 331984 62086 331996
rect 53098 331916 53104 331968
rect 53156 331956 53162 331968
rect 236242 331956 236270 331996
rect 239950 331984 239956 331996
rect 240008 331984 240014 332036
rect 294325 332027 294383 332033
rect 294325 331993 294337 332027
rect 294371 332024 294383 332027
rect 539686 332024 539692 332036
rect 294371 331996 539692 332024
rect 294371 331993 294383 331996
rect 294325 331987 294383 331993
rect 539686 331984 539692 331996
rect 539744 331984 539750 332036
rect 238018 331956 238024 331968
rect 53156 331928 236270 331956
rect 236334 331928 238024 331956
rect 53156 331916 53162 331928
rect 32398 331848 32404 331900
rect 32456 331888 32462 331900
rect 236334 331888 236362 331928
rect 238018 331916 238024 331928
rect 238076 331916 238082 331968
rect 290366 331916 290372 331968
rect 290424 331956 290430 331968
rect 538214 331956 538220 331968
rect 290424 331928 538220 331956
rect 290424 331916 290430 331928
rect 538214 331916 538220 331928
rect 538272 331916 538278 331968
rect 32456 331860 236362 331888
rect 267553 331891 267611 331897
rect 32456 331848 32462 331860
rect 267553 331857 267565 331891
rect 267599 331888 267611 331891
rect 287054 331888 287060 331900
rect 267599 331860 287060 331888
rect 267599 331857 267611 331860
rect 267553 331851 267611 331857
rect 287054 331848 287060 331860
rect 287112 331848 287118 331900
rect 295518 331848 295524 331900
rect 295576 331888 295582 331900
rect 547966 331888 547972 331900
rect 295576 331860 547972 331888
rect 295576 331848 295582 331860
rect 547966 331848 547972 331860
rect 548024 331848 548030 331900
rect 155862 331780 155868 331832
rect 155920 331820 155926 331832
rect 250714 331820 250720 331832
rect 155920 331792 250720 331820
rect 155920 331780 155926 331792
rect 250714 331780 250720 331792
rect 250772 331780 250778 331832
rect 274818 331780 274824 331832
rect 274876 331820 274882 331832
rect 385678 331820 385684 331832
rect 274876 331792 385684 331820
rect 274876 331780 274882 331792
rect 385678 331780 385684 331792
rect 385736 331780 385742 331832
rect 184842 331712 184848 331764
rect 184900 331752 184906 331764
rect 253934 331752 253940 331764
rect 184900 331724 253940 331752
rect 184900 331712 184906 331724
rect 253934 331712 253940 331724
rect 253992 331712 253998 331764
rect 271690 331712 271696 331764
rect 271748 331752 271754 331764
rect 357434 331752 357440 331764
rect 271748 331724 357440 331752
rect 271748 331712 271754 331724
rect 357434 331712 357440 331724
rect 357492 331712 357498 331764
rect 188982 331644 188988 331696
rect 189040 331684 189046 331696
rect 254302 331684 254308 331696
rect 189040 331656 254308 331684
rect 189040 331644 189046 331656
rect 254302 331644 254308 331656
rect 254360 331644 254366 331696
rect 269666 331644 269672 331696
rect 269724 331684 269730 331696
rect 338114 331684 338120 331696
rect 269724 331656 338120 331684
rect 269724 331644 269730 331656
rect 338114 331644 338120 331656
rect 338172 331644 338178 331696
rect 213822 331576 213828 331628
rect 213880 331616 213886 331628
rect 256878 331616 256884 331628
rect 213880 331588 256884 331616
rect 213880 331576 213886 331588
rect 256878 331576 256884 331588
rect 256936 331576 256942 331628
rect 276934 331576 276940 331628
rect 276992 331616 276998 331628
rect 335354 331616 335360 331628
rect 276992 331588 335360 331616
rect 276992 331576 276998 331588
rect 335354 331576 335360 331588
rect 335412 331576 335418 331628
rect 224862 331508 224868 331560
rect 224920 331548 224926 331560
rect 257982 331548 257988 331560
rect 224920 331520 257988 331548
rect 224920 331508 224926 331520
rect 257982 331508 257988 331520
rect 258040 331508 258046 331560
rect 268470 331508 268476 331560
rect 268528 331548 268534 331560
rect 324406 331548 324412 331560
rect 268528 331520 324412 331548
rect 268528 331508 268534 331520
rect 324406 331508 324412 331520
rect 324464 331508 324470 331560
rect 234338 331440 234344 331492
rect 234396 331480 234402 331492
rect 258902 331480 258908 331492
rect 234396 331452 258908 331480
rect 234396 331440 234402 331452
rect 258902 331440 258908 331452
rect 258960 331440 258966 331492
rect 267366 331440 267372 331492
rect 267424 331480 267430 331492
rect 313918 331480 313924 331492
rect 267424 331452 313924 331480
rect 267424 331440 267430 331452
rect 313918 331440 313924 331452
rect 313976 331440 313982 331492
rect 235997 331415 236055 331421
rect 235997 331381 236009 331415
rect 236043 331412 236055 331415
rect 242710 331412 242716 331424
rect 236043 331384 242716 331412
rect 236043 331381 236055 331384
rect 235997 331375 236055 331381
rect 242710 331372 242716 331384
rect 242768 331372 242774 331424
rect 266354 331372 266360 331424
rect 266412 331412 266418 331424
rect 304994 331412 305000 331424
rect 266412 331384 305000 331412
rect 266412 331372 266418 331384
rect 304994 331372 305000 331384
rect 305052 331372 305058 331424
rect 193122 331168 193128 331220
rect 193180 331208 193186 331220
rect 254670 331208 254676 331220
rect 193180 331180 254676 331208
rect 193180 331168 193186 331180
rect 254670 331168 254676 331180
rect 254728 331168 254734 331220
rect 279786 331168 279792 331220
rect 279844 331208 279850 331220
rect 434714 331208 434720 331220
rect 279844 331180 434720 331208
rect 279844 331168 279850 331180
rect 434714 331168 434720 331180
rect 434772 331168 434778 331220
rect 153010 331100 153016 331152
rect 153068 331140 153074 331152
rect 250622 331140 250628 331152
rect 153068 331112 250628 331140
rect 153068 331100 153074 331112
rect 250622 331100 250628 331112
rect 250680 331100 250686 331152
rect 293034 331100 293040 331152
rect 293092 331140 293098 331152
rect 450538 331140 450544 331152
rect 293092 331112 450544 331140
rect 293092 331100 293098 331112
rect 450538 331100 450544 331112
rect 450596 331100 450602 331152
rect 111702 331032 111708 331084
rect 111760 331072 111766 331084
rect 246574 331072 246580 331084
rect 111760 331044 246580 331072
rect 111760 331032 111766 331044
rect 246574 331032 246580 331044
rect 246632 331032 246638 331084
rect 285306 331032 285312 331084
rect 285364 331072 285370 331084
rect 488534 331072 488540 331084
rect 285364 331044 488540 331072
rect 285364 331032 285370 331044
rect 488534 331032 488540 331044
rect 488592 331032 488598 331084
rect 108942 330964 108948 331016
rect 109000 331004 109006 331016
rect 245746 331004 245752 331016
rect 109000 330976 245752 331004
rect 109000 330964 109006 330976
rect 245746 330964 245752 330976
rect 245804 330964 245810 331016
rect 284294 331004 284300 331016
rect 273226 330976 284300 331004
rect 102042 330896 102048 330948
rect 102100 330936 102106 330948
rect 245286 330936 245292 330948
rect 102100 330908 245292 330936
rect 102100 330896 102106 330908
rect 245286 330896 245292 330908
rect 245344 330896 245350 330948
rect 79318 330828 79324 330880
rect 79376 330868 79382 330880
rect 242802 330868 242808 330880
rect 79376 330840 242808 330868
rect 79376 330828 79382 330840
rect 242802 330828 242808 330840
rect 242860 330828 242866 330880
rect 264241 330871 264299 330877
rect 264241 330837 264253 330871
rect 264287 330868 264299 330871
rect 273226 330868 273254 330976
rect 284294 330964 284300 330976
rect 284352 330964 284358 331016
rect 285582 330964 285588 331016
rect 285640 331004 285646 331016
rect 490558 331004 490564 331016
rect 285640 330976 490564 331004
rect 285640 330964 285646 330976
rect 490558 330964 490564 330976
rect 490616 330964 490622 331016
rect 286686 330896 286692 330948
rect 286744 330936 286750 330948
rect 502334 330936 502340 330948
rect 286744 330908 502340 330936
rect 286744 330896 286750 330908
rect 502334 330896 502340 330908
rect 502392 330896 502398 330948
rect 264287 330840 273254 330868
rect 264287 330837 264299 330840
rect 264241 330831 264299 330837
rect 287790 330828 287796 330880
rect 287848 330868 287854 330880
rect 512638 330868 512644 330880
rect 287848 330840 512644 330868
rect 287848 330828 287854 330840
rect 512638 330828 512644 330840
rect 512696 330828 512702 330880
rect 68278 330760 68284 330812
rect 68336 330800 68342 330812
rect 241790 330800 241796 330812
rect 68336 330772 241796 330800
rect 68336 330760 68342 330772
rect 241790 330760 241796 330772
rect 241848 330760 241854 330812
rect 272886 330760 272892 330812
rect 272944 330760 272950 330812
rect 299934 330760 299940 330812
rect 299992 330800 299998 330812
rect 536834 330800 536840 330812
rect 299992 330772 536840 330800
rect 299992 330760 299998 330772
rect 536834 330760 536840 330772
rect 536892 330760 536898 330812
rect 57238 330692 57244 330744
rect 57296 330732 57302 330744
rect 240318 330732 240324 330744
rect 57296 330704 240324 330732
rect 57296 330692 57302 330704
rect 240318 330692 240324 330704
rect 240376 330692 240382 330744
rect 39298 330624 39304 330676
rect 39356 330664 39362 330676
rect 238938 330664 238944 330676
rect 39356 330636 238944 330664
rect 39356 330624 39362 330636
rect 238938 330624 238944 330636
rect 238996 330624 239002 330676
rect 37182 330556 37188 330608
rect 37240 330596 37246 330608
rect 230293 330599 230351 330605
rect 230293 330596 230305 330599
rect 37240 330568 230305 330596
rect 37240 330556 37246 330568
rect 230293 330565 230305 330568
rect 230339 330565 230351 330599
rect 236270 330596 236276 330608
rect 230293 330559 230351 330565
rect 230400 330568 236276 330596
rect 22738 330488 22744 330540
rect 22796 330528 22802 330540
rect 230400 330528 230428 330568
rect 236270 330556 236276 330568
rect 236328 330556 236334 330608
rect 22796 330500 230428 330528
rect 22796 330488 22802 330500
rect 255590 330488 255596 330540
rect 255648 330528 255654 330540
rect 256234 330528 256240 330540
rect 255648 330500 256240 330528
rect 255648 330488 255654 330500
rect 256234 330488 256240 330500
rect 256292 330488 256298 330540
rect 258626 330488 258632 330540
rect 258684 330528 258690 330540
rect 259270 330528 259276 330540
rect 258684 330500 259276 330528
rect 258684 330488 258690 330500
rect 259270 330488 259276 330500
rect 259328 330488 259334 330540
rect 267182 330488 267188 330540
rect 267240 330528 267246 330540
rect 267458 330528 267464 330540
rect 267240 330500 267464 330528
rect 267240 330488 267246 330500
rect 267458 330488 267464 330500
rect 267516 330488 267522 330540
rect 195882 330420 195888 330472
rect 195940 330460 195946 330472
rect 255038 330460 255044 330472
rect 195940 330432 255044 330460
rect 195940 330420 195946 330432
rect 255038 330420 255044 330432
rect 255096 330420 255102 330472
rect 255406 330420 255412 330472
rect 255464 330460 255470 330472
rect 255958 330460 255964 330472
rect 255464 330432 255964 330460
rect 255464 330420 255470 330432
rect 255958 330420 255964 330432
rect 256016 330420 256022 330472
rect 259638 330420 259644 330472
rect 259696 330460 259702 330472
rect 260282 330460 260288 330472
rect 259696 330432 260288 330460
rect 259696 330420 259702 330432
rect 260282 330420 260288 330432
rect 260340 330420 260346 330472
rect 272150 330420 272156 330472
rect 272208 330460 272214 330472
rect 272794 330460 272800 330472
rect 272208 330432 272800 330460
rect 272208 330420 272214 330432
rect 272794 330420 272800 330432
rect 272852 330420 272858 330472
rect 272904 330460 272932 330760
rect 289262 330692 289268 330744
rect 289320 330732 289326 330744
rect 528646 330732 528652 330744
rect 289320 330704 528652 330732
rect 289320 330692 289326 330704
rect 528646 330692 528652 330704
rect 528704 330692 528710 330744
rect 291102 330624 291108 330676
rect 291160 330664 291166 330676
rect 546494 330664 546500 330676
rect 291160 330636 546500 330664
rect 291160 330624 291166 330636
rect 546494 330624 546500 330636
rect 546552 330624 546558 330676
rect 293310 330556 293316 330608
rect 293368 330596 293374 330608
rect 293368 330568 295104 330596
rect 293368 330556 293374 330568
rect 294046 330488 294052 330540
rect 294104 330528 294110 330540
rect 294782 330528 294788 330540
rect 294104 330500 294788 330528
rect 294104 330488 294110 330500
rect 294782 330488 294788 330500
rect 294840 330488 294846 330540
rect 295076 330528 295104 330568
rect 295794 330556 295800 330608
rect 295852 330596 295858 330608
rect 564526 330596 564532 330608
rect 295852 330568 564532 330596
rect 295852 330556 295858 330568
rect 564526 330556 564532 330568
rect 564584 330556 564590 330608
rect 565814 330528 565820 330540
rect 295076 330500 565820 330528
rect 565814 330488 565820 330500
rect 565872 330488 565878 330540
rect 273070 330460 273076 330472
rect 272904 330432 273076 330460
rect 273070 330420 273076 330432
rect 273128 330420 273134 330472
rect 274082 330420 274088 330472
rect 274140 330460 274146 330472
rect 375374 330460 375380 330472
rect 274140 330432 375380 330460
rect 274140 330420 274146 330432
rect 375374 330420 375380 330432
rect 375432 330420 375438 330472
rect 202782 330352 202788 330404
rect 202840 330392 202846 330404
rect 254854 330392 254860 330404
rect 202840 330364 254860 330392
rect 202840 330352 202846 330364
rect 254854 330352 254860 330364
rect 254912 330352 254918 330404
rect 257246 330392 257252 330404
rect 254964 330364 257252 330392
rect 217962 330284 217968 330336
rect 218020 330324 218026 330336
rect 254964 330324 254992 330364
rect 257246 330352 257252 330364
rect 257304 330352 257310 330404
rect 270402 330352 270408 330404
rect 270460 330392 270466 330404
rect 342898 330392 342904 330404
rect 270460 330364 342904 330392
rect 270460 330352 270466 330364
rect 342898 330352 342904 330364
rect 342956 330352 342962 330404
rect 255774 330324 255780 330336
rect 218020 330296 254992 330324
rect 255735 330296 255780 330324
rect 218020 330284 218026 330296
rect 255774 330284 255780 330296
rect 255832 330284 255838 330336
rect 255866 330284 255872 330336
rect 255924 330324 255930 330336
rect 256326 330324 256332 330336
rect 255924 330296 256332 330324
rect 255924 330284 255930 330296
rect 256326 330284 256332 330296
rect 256384 330284 256390 330336
rect 260834 330284 260840 330336
rect 260892 330324 260898 330336
rect 261110 330324 261116 330336
rect 260892 330296 261116 330324
rect 260892 330284 260898 330296
rect 261110 330284 261116 330296
rect 261168 330284 261174 330336
rect 268930 330284 268936 330336
rect 268988 330324 268994 330336
rect 328454 330324 328460 330336
rect 268988 330296 328460 330324
rect 268988 330284 268994 330296
rect 328454 330284 328460 330296
rect 328512 330284 328518 330336
rect 220722 330216 220728 330268
rect 220780 330256 220786 330268
rect 220780 330228 244274 330256
rect 220780 330216 220786 330228
rect 230293 330191 230351 330197
rect 230293 330157 230305 330191
rect 230339 330188 230351 330191
rect 238570 330188 238576 330200
rect 230339 330160 238576 330188
rect 230339 330157 230351 330160
rect 230293 330151 230351 330157
rect 238570 330148 238576 330160
rect 238628 330148 238634 330200
rect 244246 330188 244274 330228
rect 255406 330216 255412 330268
rect 255464 330256 255470 330268
rect 256602 330256 256608 330268
rect 255464 330228 256608 330256
rect 255464 330216 255470 330228
rect 256602 330216 256608 330228
rect 256660 330216 256666 330268
rect 267642 330216 267648 330268
rect 267700 330256 267706 330268
rect 317414 330256 317420 330268
rect 267700 330228 317420 330256
rect 267700 330216 267706 330228
rect 317414 330216 317420 330228
rect 317472 330216 317478 330268
rect 257614 330188 257620 330200
rect 244246 330160 257620 330188
rect 257614 330148 257620 330160
rect 257672 330148 257678 330200
rect 261110 330148 261116 330200
rect 261168 330188 261174 330200
rect 261570 330188 261576 330200
rect 261168 330160 261576 330188
rect 261168 330148 261174 330160
rect 261570 330148 261576 330160
rect 261628 330148 261634 330200
rect 263870 330148 263876 330200
rect 263928 330188 263934 330200
rect 264238 330188 264244 330200
rect 263928 330160 264244 330188
rect 263928 330148 263934 330160
rect 264238 330148 264244 330160
rect 264296 330148 264302 330200
rect 275094 329740 275100 329792
rect 275152 329780 275158 329792
rect 389818 329780 389824 329792
rect 275152 329752 389824 329780
rect 275152 329740 275158 329752
rect 389818 329740 389824 329752
rect 389876 329740 389882 329792
rect 146202 329672 146208 329724
rect 146260 329712 146266 329724
rect 249978 329712 249984 329724
rect 146260 329684 249984 329712
rect 146260 329672 146266 329684
rect 249978 329672 249984 329684
rect 250036 329672 250042 329724
rect 276842 329672 276848 329724
rect 276900 329712 276906 329724
rect 407114 329712 407120 329724
rect 276900 329684 407120 329712
rect 276900 329672 276906 329684
rect 407114 329672 407120 329684
rect 407172 329672 407178 329724
rect 99282 329604 99288 329656
rect 99340 329644 99346 329656
rect 245013 329647 245071 329653
rect 245013 329644 245025 329647
rect 99340 329616 245025 329644
rect 99340 329604 99346 329616
rect 245013 329613 245025 329616
rect 245059 329613 245071 329647
rect 245013 329607 245071 329613
rect 277210 329604 277216 329656
rect 277268 329644 277274 329656
rect 409874 329644 409880 329656
rect 277268 329616 409880 329644
rect 277268 329604 277274 329616
rect 409874 329604 409880 329616
rect 409932 329604 409938 329656
rect 93118 329536 93124 329588
rect 93176 329576 93182 329588
rect 244366 329576 244372 329588
rect 93176 329548 244372 329576
rect 93176 329536 93182 329548
rect 244366 329536 244372 329548
rect 244424 329536 244430 329588
rect 280062 329536 280068 329588
rect 280120 329576 280126 329588
rect 438854 329576 438860 329588
rect 280120 329548 438860 329576
rect 280120 329536 280126 329548
rect 438854 329536 438860 329548
rect 438912 329536 438918 329588
rect 75178 329468 75184 329520
rect 75236 329508 75242 329520
rect 242526 329508 242532 329520
rect 75236 329480 242532 329508
rect 75236 329468 75242 329480
rect 242526 329468 242532 329480
rect 242584 329468 242590 329520
rect 283650 329468 283656 329520
rect 283708 329508 283714 329520
rect 474734 329508 474740 329520
rect 283708 329480 474740 329508
rect 283708 329468 283714 329480
rect 474734 329468 474740 329480
rect 474792 329468 474798 329520
rect 71038 329400 71044 329452
rect 71096 329440 71102 329452
rect 242158 329440 242164 329452
rect 71096 329412 242164 329440
rect 71096 329400 71102 329412
rect 242158 329400 242164 329412
rect 242216 329400 242222 329452
rect 288250 329400 288256 329452
rect 288308 329440 288314 329452
rect 517514 329440 517520 329452
rect 288308 329412 517520 329440
rect 288308 329400 288314 329412
rect 517514 329400 517520 329412
rect 517572 329400 517578 329452
rect 63402 329332 63408 329384
rect 63460 329372 63466 329384
rect 241422 329372 241428 329384
rect 63460 329344 241428 329372
rect 63460 329332 63466 329344
rect 241422 329332 241428 329344
rect 241480 329332 241486 329384
rect 289630 329332 289636 329384
rect 289688 329372 289694 329384
rect 530578 329372 530584 329384
rect 289688 329344 530584 329372
rect 289688 329332 289694 329344
rect 530578 329332 530584 329344
rect 530636 329332 530642 329384
rect 61378 329264 61384 329316
rect 61436 329304 61442 329316
rect 241054 329304 241060 329316
rect 61436 329276 241060 329304
rect 61436 329264 61442 329276
rect 241054 329264 241060 329276
rect 241112 329264 241118 329316
rect 304166 329264 304172 329316
rect 304224 329304 304230 329316
rect 561674 329304 561680 329316
rect 304224 329276 561680 329304
rect 304224 329264 304230 329276
rect 561674 329264 561680 329276
rect 561732 329264 561738 329316
rect 57330 329196 57336 329248
rect 57388 329236 57394 329248
rect 240686 329236 240692 329248
rect 57388 329208 240692 329236
rect 57388 329196 57394 329208
rect 240686 329196 240692 329208
rect 240744 329196 240750 329248
rect 291838 329196 291844 329248
rect 291896 329236 291902 329248
rect 551278 329236 551284 329248
rect 291896 329208 551284 329236
rect 291896 329196 291902 329208
rect 551278 329196 551284 329208
rect 551336 329196 551342 329248
rect 39390 329128 39396 329180
rect 39448 329168 39454 329180
rect 236822 329168 236828 329180
rect 39448 329140 236828 329168
rect 39448 329128 39454 329140
rect 236822 329128 236828 329140
rect 236880 329128 236886 329180
rect 291746 329128 291752 329180
rect 291804 329168 291810 329180
rect 556154 329168 556160 329180
rect 291804 329140 556160 329168
rect 291804 329128 291810 329140
rect 556154 329128 556160 329140
rect 556212 329128 556218 329180
rect 32490 329060 32496 329112
rect 32548 329100 32554 329112
rect 238110 329100 238116 329112
rect 32548 329072 238116 329100
rect 32548 329060 32554 329072
rect 238110 329060 238116 329072
rect 238168 329060 238174 329112
rect 264882 329060 264888 329112
rect 264940 329100 264946 329112
rect 291194 329100 291200 329112
rect 264940 329072 291200 329100
rect 264940 329060 264946 329072
rect 291194 329060 291200 329072
rect 291252 329060 291258 329112
rect 294233 329103 294291 329109
rect 294233 329069 294245 329103
rect 294279 329100 294291 329103
rect 569954 329100 569960 329112
rect 294279 329072 569960 329100
rect 294279 329069 294291 329072
rect 294233 329063 294291 329069
rect 569954 329060 569960 329072
rect 570012 329060 570018 329112
rect 273622 328992 273628 329044
rect 273680 329032 273686 329044
rect 378778 329032 378784 329044
rect 273680 329004 378784 329032
rect 273680 328992 273686 329004
rect 378778 328992 378784 329004
rect 378836 328992 378842 329044
rect 270034 328924 270040 328976
rect 270092 328964 270098 328976
rect 340874 328964 340880 328976
rect 270092 328936 340880 328964
rect 270092 328924 270098 328936
rect 340874 328924 340880 328936
rect 340932 328924 340938 328976
rect 270126 328692 270132 328704
rect 270087 328664 270132 328692
rect 270126 328652 270132 328664
rect 270184 328652 270190 328704
rect 273438 328380 273444 328432
rect 273496 328420 273502 328432
rect 382274 328420 382280 328432
rect 273496 328392 382280 328420
rect 273496 328380 273502 328392
rect 382274 328380 382280 328392
rect 382332 328380 382338 328432
rect 275738 328312 275744 328364
rect 275796 328352 275802 328364
rect 392578 328352 392584 328364
rect 275796 328324 392584 328352
rect 275796 328312 275802 328324
rect 392578 328312 392584 328324
rect 392636 328312 392642 328364
rect 265894 328244 265900 328296
rect 265952 328284 265958 328296
rect 266170 328284 266176 328296
rect 265952 328256 266176 328284
rect 265952 328244 265958 328256
rect 266170 328244 266176 328256
rect 266228 328244 266234 328296
rect 278314 328244 278320 328296
rect 278372 328284 278378 328296
rect 414014 328284 414020 328296
rect 278372 328256 414020 328284
rect 278372 328244 278378 328256
rect 414014 328244 414020 328256
rect 414072 328244 414078 328296
rect 119982 328176 119988 328228
rect 120040 328216 120046 328228
rect 245102 328216 245108 328228
rect 120040 328188 245108 328216
rect 120040 328176 120046 328188
rect 245102 328176 245108 328188
rect 245160 328176 245166 328228
rect 277854 328176 277860 328228
rect 277912 328216 277918 328228
rect 416774 328216 416780 328228
rect 277912 328188 416780 328216
rect 277912 328176 277918 328188
rect 416774 328176 416780 328188
rect 416832 328176 416838 328228
rect 113082 328108 113088 328160
rect 113140 328148 113146 328160
rect 246390 328148 246396 328160
rect 113140 328120 246396 328148
rect 113140 328108 113146 328120
rect 246390 328108 246396 328120
rect 246448 328108 246454 328160
rect 278222 328108 278228 328160
rect 278280 328148 278286 328160
rect 420914 328148 420920 328160
rect 278280 328120 420920 328148
rect 278280 328108 278286 328120
rect 420914 328108 420920 328120
rect 420972 328108 420978 328160
rect 111058 328040 111064 328092
rect 111116 328080 111122 328092
rect 246022 328080 246028 328092
rect 111116 328052 246028 328080
rect 111116 328040 111122 328052
rect 246022 328040 246028 328052
rect 246080 328040 246086 328092
rect 293678 328040 293684 328092
rect 293736 328080 293742 328092
rect 453298 328080 453304 328092
rect 293736 328052 453304 328080
rect 293736 328040 293742 328052
rect 453298 328040 453304 328052
rect 453356 328040 453362 328092
rect 106182 327972 106188 328024
rect 106240 328012 106246 328024
rect 245838 328012 245844 328024
rect 106240 327984 245844 328012
rect 106240 327972 106246 327984
rect 245838 327972 245844 327984
rect 245896 327972 245902 328024
rect 290918 327972 290924 328024
rect 290976 328012 290982 328024
rect 464338 328012 464344 328024
rect 290976 327984 464344 328012
rect 290976 327972 290982 327984
rect 464338 327972 464344 327984
rect 464396 327972 464402 328024
rect 95050 327904 95056 327956
rect 95108 327944 95114 327956
rect 244734 327944 244740 327956
rect 95108 327916 244740 327944
rect 95108 327904 95114 327916
rect 244734 327904 244740 327916
rect 244792 327904 244798 327956
rect 286502 327904 286508 327956
rect 286560 327944 286566 327956
rect 466454 327944 466460 327956
rect 286560 327916 466460 327944
rect 286560 327904 286566 327916
rect 466454 327904 466460 327916
rect 466512 327904 466518 327956
rect 43438 327836 43444 327888
rect 43496 327876 43502 327888
rect 237282 327876 237288 327888
rect 43496 327848 237288 327876
rect 43496 327836 43502 327848
rect 237282 327836 237288 327848
rect 237340 327836 237346 327888
rect 284110 327836 284116 327888
rect 284168 327876 284174 327888
rect 477494 327876 477500 327888
rect 284168 327848 477500 327876
rect 284168 327836 284174 327848
rect 477494 327836 477500 327848
rect 477552 327836 477558 327888
rect 45462 327768 45468 327820
rect 45520 327808 45526 327820
rect 239306 327808 239312 327820
rect 45520 327780 239312 327808
rect 45520 327768 45526 327780
rect 239306 327768 239312 327780
rect 239364 327768 239370 327820
rect 286778 327768 286784 327820
rect 286836 327808 286842 327820
rect 503714 327808 503720 327820
rect 286836 327780 503720 327808
rect 286836 327768 286842 327780
rect 503714 327768 503720 327780
rect 503772 327768 503778 327820
rect 28902 327700 28908 327752
rect 28960 327740 28966 327752
rect 237466 327740 237472 327752
rect 28960 327712 237472 327740
rect 28960 327700 28966 327712
rect 237466 327700 237472 327712
rect 237524 327700 237530 327752
rect 292114 327700 292120 327752
rect 292172 327740 292178 327752
rect 560294 327740 560300 327752
rect 292172 327712 560300 327740
rect 292172 327700 292178 327712
rect 560294 327700 560300 327712
rect 560352 327700 560358 327752
rect 275554 326884 275560 326936
rect 275612 326924 275618 326936
rect 396718 326924 396724 326936
rect 275612 326896 396724 326924
rect 275612 326884 275618 326896
rect 396718 326884 396724 326896
rect 396776 326884 396782 326936
rect 278590 326816 278596 326868
rect 278648 326856 278654 326868
rect 423766 326856 423772 326868
rect 278648 326828 423772 326856
rect 278648 326816 278654 326828
rect 423766 326816 423772 326828
rect 423824 326816 423830 326868
rect 285398 326748 285404 326800
rect 285456 326788 285462 326800
rect 290645 326791 290703 326797
rect 290645 326788 290657 326791
rect 285456 326760 290657 326788
rect 285456 326748 285462 326760
rect 290645 326757 290657 326760
rect 290691 326757 290703 326791
rect 290645 326751 290703 326757
rect 293586 326748 293592 326800
rect 293644 326788 293650 326800
rect 443638 326788 443644 326800
rect 293644 326760 443644 326788
rect 293644 326748 293650 326760
rect 443638 326748 443644 326760
rect 443696 326748 443702 326800
rect 234982 326720 234988 326732
rect 234943 326692 234988 326720
rect 234982 326680 234988 326692
rect 235040 326680 235046 326732
rect 235813 326723 235871 326729
rect 235813 326689 235825 326723
rect 235859 326720 235871 326723
rect 241606 326720 241612 326732
rect 235859 326692 241612 326720
rect 235859 326689 235871 326692
rect 235813 326683 235871 326689
rect 241606 326680 241612 326692
rect 241664 326680 241670 326732
rect 284938 326680 284944 326732
rect 284996 326720 285002 326732
rect 284996 326692 290504 326720
rect 284996 326680 285002 326692
rect 117222 326612 117228 326664
rect 117280 326652 117286 326664
rect 246850 326652 246856 326664
rect 117280 326624 246856 326652
rect 117280 326612 117286 326624
rect 246850 326612 246856 326624
rect 246908 326612 246914 326664
rect 68370 326544 68376 326596
rect 68428 326584 68434 326596
rect 235813 326587 235871 326593
rect 235813 326584 235825 326587
rect 68428 326556 235825 326584
rect 68428 326544 68434 326556
rect 235813 326553 235825 326556
rect 235859 326553 235871 326587
rect 240870 326584 240876 326596
rect 235813 326547 235871 326553
rect 235920 326556 240876 326584
rect 58618 326476 58624 326528
rect 58676 326516 58682 326528
rect 235920 326516 235948 326556
rect 240870 326544 240876 326556
rect 240928 326544 240934 326596
rect 280614 326584 280620 326596
rect 280575 326556 280620 326584
rect 280614 326544 280620 326556
rect 280672 326544 280678 326596
rect 286870 326544 286876 326596
rect 286928 326584 286934 326596
rect 290476 326584 290504 326692
rect 290550 326680 290556 326732
rect 290608 326720 290614 326732
rect 461578 326720 461584 326732
rect 290608 326692 461584 326720
rect 290608 326680 290614 326692
rect 461578 326680 461584 326692
rect 461636 326680 461642 326732
rect 290645 326655 290703 326661
rect 290645 326621 290657 326655
rect 290691 326652 290703 326655
rect 481726 326652 481732 326664
rect 290691 326624 481732 326652
rect 290691 326621 290703 326624
rect 290645 326615 290703 326621
rect 481726 326612 481732 326624
rect 481784 326612 481790 326664
rect 485774 326584 485780 326596
rect 286928 326556 290412 326584
rect 290476 326556 485780 326584
rect 286928 326544 286934 326556
rect 240042 326516 240048 326528
rect 58676 326488 235948 326516
rect 236012 326488 240048 326516
rect 58676 326476 58682 326488
rect 50982 326408 50988 326460
rect 51040 326448 51046 326460
rect 236012 326448 236040 326488
rect 240042 326476 240048 326488
rect 240100 326476 240106 326528
rect 288066 326476 288072 326528
rect 288124 326516 288130 326528
rect 290384 326516 290412 326556
rect 485774 326544 485780 326556
rect 485832 326544 485838 326596
rect 492674 326516 492680 326528
rect 288124 326488 290320 326516
rect 290384 326488 492680 326516
rect 288124 326476 288130 326488
rect 238478 326448 238484 326460
rect 51040 326420 236040 326448
rect 236104 326420 238484 326448
rect 51040 326408 51046 326420
rect 35802 326340 35808 326392
rect 35860 326380 35866 326392
rect 236104 326380 236132 326420
rect 238478 326408 238484 326420
rect 238536 326408 238542 326460
rect 243078 326408 243084 326460
rect 243136 326448 243142 326460
rect 244090 326448 244096 326460
rect 243136 326420 244096 326448
rect 243136 326408 243142 326420
rect 244090 326408 244096 326420
rect 244148 326408 244154 326460
rect 273806 326408 273812 326460
rect 273864 326448 273870 326460
rect 274542 326448 274548 326460
rect 273864 326420 274548 326448
rect 273864 326408 273870 326420
rect 274542 326408 274548 326420
rect 274600 326408 274606 326460
rect 281350 326408 281356 326460
rect 281408 326408 281414 326460
rect 282362 326408 282368 326460
rect 282420 326448 282426 326460
rect 282546 326448 282552 326460
rect 282420 326420 282552 326448
rect 282420 326408 282426 326420
rect 282546 326408 282552 326420
rect 282604 326408 282610 326460
rect 289446 326408 289452 326460
rect 289504 326448 289510 326460
rect 290292 326448 290320 326488
rect 492674 326476 492680 326488
rect 492732 326476 492738 326528
rect 506566 326448 506572 326460
rect 289504 326420 289860 326448
rect 290292 326420 506572 326448
rect 289504 326408 289510 326420
rect 35860 326352 236132 326380
rect 35860 326340 35866 326352
rect 236178 326340 236184 326392
rect 236236 326380 236242 326392
rect 236546 326380 236552 326392
rect 236236 326352 236552 326380
rect 236236 326340 236242 326352
rect 236546 326340 236552 326352
rect 236604 326340 236610 326392
rect 237374 326340 237380 326392
rect 237432 326380 237438 326392
rect 237926 326380 237932 326392
rect 237432 326352 237932 326380
rect 237432 326340 237438 326352
rect 237926 326340 237932 326352
rect 237984 326340 237990 326392
rect 239030 326340 239036 326392
rect 239088 326380 239094 326392
rect 239398 326380 239404 326392
rect 239088 326352 239404 326380
rect 239088 326340 239094 326352
rect 239398 326340 239404 326352
rect 239456 326340 239462 326392
rect 243170 326340 243176 326392
rect 243228 326380 243234 326392
rect 243722 326380 243728 326392
rect 243228 326352 243728 326380
rect 243228 326340 243234 326352
rect 243722 326340 243728 326352
rect 243780 326340 243786 326392
rect 246114 326340 246120 326392
rect 246172 326380 246178 326392
rect 246942 326380 246948 326392
rect 246172 326352 246948 326380
rect 246172 326340 246178 326352
rect 246942 326340 246948 326352
rect 247000 326340 247006 326392
rect 247126 326340 247132 326392
rect 247184 326380 247190 326392
rect 248230 326380 248236 326392
rect 247184 326352 248236 326380
rect 247184 326340 247190 326352
rect 248230 326340 248236 326352
rect 248288 326340 248294 326392
rect 248690 326340 248696 326392
rect 248748 326380 248754 326392
rect 249150 326380 249156 326392
rect 248748 326352 249156 326380
rect 248748 326340 248754 326352
rect 249150 326340 249156 326352
rect 249208 326340 249214 326392
rect 273530 326340 273536 326392
rect 273588 326380 273594 326392
rect 273990 326380 273996 326392
rect 273588 326352 273996 326380
rect 273588 326340 273594 326352
rect 273990 326340 273996 326352
rect 274048 326340 274054 326392
rect 275002 326340 275008 326392
rect 275060 326380 275066 326392
rect 275370 326380 275376 326392
rect 275060 326352 275376 326380
rect 275060 326340 275066 326352
rect 275370 326340 275376 326352
rect 275428 326340 275434 326392
rect 280338 326340 280344 326392
rect 280396 326380 280402 326392
rect 280982 326380 280988 326392
rect 280396 326352 280988 326380
rect 280396 326340 280402 326352
rect 280982 326340 280988 326352
rect 281040 326340 281046 326392
rect 280614 326312 280620 326324
rect 280575 326284 280620 326312
rect 280614 326272 280620 326284
rect 280672 326272 280678 326324
rect 235166 326204 235172 326256
rect 235224 326244 235230 326256
rect 235626 326244 235632 326256
rect 235224 326216 235632 326244
rect 235224 326204 235230 326216
rect 235626 326204 235632 326216
rect 235684 326204 235690 326256
rect 247218 326204 247224 326256
rect 247276 326244 247282 326256
rect 247402 326244 247408 326256
rect 247276 326216 247408 326244
rect 247276 326204 247282 326216
rect 247402 326204 247408 326216
rect 247460 326204 247466 326256
rect 247494 326204 247500 326256
rect 247552 326244 247558 326256
rect 247678 326244 247684 326256
rect 247552 326216 247684 326244
rect 247552 326204 247558 326216
rect 247678 326204 247684 326216
rect 247736 326204 247742 326256
rect 281368 326244 281396 326408
rect 288986 326340 288992 326392
rect 289044 326380 289050 326392
rect 289722 326380 289728 326392
rect 289044 326352 289728 326380
rect 289044 326340 289050 326352
rect 289722 326340 289728 326352
rect 289780 326340 289786 326392
rect 289832 326380 289860 326420
rect 506566 326408 506572 326420
rect 506624 326408 506630 326460
rect 519538 326380 519544 326392
rect 289832 326352 519544 326380
rect 519538 326340 519544 326352
rect 519596 326340 519602 326392
rect 281442 326244 281448 326256
rect 281368 326216 281448 326244
rect 281442 326204 281448 326216
rect 281500 326204 281506 326256
rect 282270 326204 282276 326256
rect 282328 326244 282334 326256
rect 282638 326244 282644 326256
rect 282328 326216 282644 326244
rect 282328 326204 282334 326216
rect 282638 326204 282644 326216
rect 282696 326204 282702 326256
rect 281718 326136 281724 326188
rect 281776 326176 281782 326188
rect 282822 326176 282828 326188
rect 281776 326148 282828 326176
rect 281776 326136 281782 326148
rect 282822 326136 282828 326148
rect 282880 326136 282886 326188
rect 247218 326068 247224 326120
rect 247276 326108 247282 326120
rect 248322 326108 248328 326120
rect 247276 326080 248328 326108
rect 247276 326068 247282 326080
rect 248322 326068 248328 326080
rect 248380 326068 248386 326120
rect 281810 326068 281816 326120
rect 281868 326108 281874 326120
rect 282270 326108 282276 326120
rect 281868 326080 282276 326108
rect 281868 326068 281874 326080
rect 282270 326068 282276 326080
rect 282328 326068 282334 326120
rect 309778 325592 309784 325644
rect 309836 325632 309842 325644
rect 580166 325632 580172 325644
rect 309836 325604 580172 325632
rect 309836 325592 309842 325604
rect 580166 325592 580172 325604
rect 580224 325592 580230 325644
rect 266630 325388 266636 325440
rect 266688 325428 266694 325440
rect 311894 325428 311900 325440
rect 266688 325400 311900 325428
rect 266688 325388 266694 325400
rect 311894 325388 311900 325400
rect 311952 325388 311958 325440
rect 268746 325320 268752 325372
rect 268804 325360 268810 325372
rect 322934 325360 322940 325372
rect 268804 325332 322940 325360
rect 268804 325320 268810 325332
rect 322934 325320 322940 325332
rect 322992 325320 322998 325372
rect 276290 325252 276296 325304
rect 276348 325292 276354 325304
rect 400214 325292 400220 325304
rect 276348 325264 400220 325292
rect 276348 325252 276354 325264
rect 400214 325252 400220 325264
rect 400272 325252 400278 325304
rect 292298 325184 292304 325236
rect 292356 325224 292362 325236
rect 457438 325224 457444 325236
rect 292356 325196 457444 325224
rect 292356 325184 292362 325196
rect 457438 325184 457444 325196
rect 457496 325184 457502 325236
rect 115198 325116 115204 325168
rect 115256 325156 115262 325168
rect 242250 325156 242256 325168
rect 115256 325128 242256 325156
rect 115256 325116 115262 325128
rect 242250 325116 242256 325128
rect 242308 325116 242314 325168
rect 286042 325116 286048 325168
rect 286100 325156 286106 325168
rect 496814 325156 496820 325168
rect 286100 325128 496820 325156
rect 286100 325116 286106 325128
rect 496814 325116 496820 325128
rect 496872 325116 496878 325168
rect 107562 325048 107568 325100
rect 107620 325088 107626 325100
rect 245930 325088 245936 325100
rect 107620 325060 245936 325088
rect 107620 325048 107626 325060
rect 245930 325048 245936 325060
rect 245988 325048 245994 325100
rect 252922 325048 252928 325100
rect 252980 325088 252986 325100
rect 252980 325060 253060 325088
rect 252980 325048 252986 325060
rect 69658 324980 69664 325032
rect 69716 325020 69722 325032
rect 242066 325020 242072 325032
rect 69716 324992 242072 325020
rect 69716 324980 69722 324992
rect 242066 324980 242072 324992
rect 242124 324980 242130 325032
rect 53742 324912 53748 324964
rect 53800 324952 53806 324964
rect 240502 324952 240508 324964
rect 53800 324924 240508 324952
rect 53800 324912 53806 324924
rect 240502 324912 240508 324924
rect 240560 324912 240566 324964
rect 253032 324896 253060 325060
rect 288158 325048 288164 325100
rect 288216 325088 288222 325100
rect 510614 325088 510620 325100
rect 288216 325060 510620 325088
rect 288216 325048 288222 325060
rect 510614 325048 510620 325060
rect 510672 325048 510678 325100
rect 289538 324980 289544 325032
rect 289596 325020 289602 325032
rect 524414 325020 524420 325032
rect 289596 324992 524420 325020
rect 289596 324980 289602 324992
rect 524414 324980 524420 324992
rect 524472 324980 524478 325032
rect 290826 324912 290832 324964
rect 290884 324952 290890 324964
rect 542354 324952 542360 324964
rect 290884 324924 542360 324952
rect 290884 324912 290890 324924
rect 542354 324912 542360 324924
rect 542412 324912 542418 324964
rect 253014 324844 253020 324896
rect 253072 324844 253078 324896
rect 268838 323892 268844 323944
rect 268896 323932 268902 323944
rect 329834 323932 329840 323944
rect 268896 323904 329840 323932
rect 268896 323892 268902 323904
rect 329834 323892 329840 323904
rect 329892 323892 329898 323944
rect 276658 323824 276664 323876
rect 276716 323864 276722 323876
rect 403618 323864 403624 323876
rect 276716 323836 403624 323864
rect 276716 323824 276722 323836
rect 403618 323824 403624 323836
rect 403676 323824 403682 323876
rect 293402 323756 293408 323808
rect 293460 323796 293466 323808
rect 447778 323796 447784 323808
rect 293460 323768 447784 323796
rect 293460 323756 293466 323768
rect 447778 323756 447784 323768
rect 447836 323756 447842 323808
rect 291562 323688 291568 323740
rect 291620 323728 291626 323740
rect 454678 323728 454684 323740
rect 291620 323700 454684 323728
rect 291620 323688 291626 323700
rect 454678 323688 454684 323700
rect 454736 323688 454742 323740
rect 286410 323620 286416 323672
rect 286468 323660 286474 323672
rect 499574 323660 499580 323672
rect 286468 323632 499580 323660
rect 286468 323620 286474 323632
rect 499574 323620 499580 323632
rect 499632 323620 499638 323672
rect 234982 323592 234988 323604
rect 234943 323564 234988 323592
rect 234982 323552 234988 323564
rect 235040 323552 235046 323604
rect 287238 323552 287244 323604
rect 287296 323592 287302 323604
rect 514846 323592 514852 323604
rect 287296 323564 514852 323592
rect 287296 323552 287302 323564
rect 514846 323552 514852 323564
rect 514904 323552 514910 323604
rect 251358 323008 251364 323060
rect 251416 323048 251422 323060
rect 251726 323048 251732 323060
rect 251416 323020 251732 323048
rect 251416 323008 251422 323020
rect 251726 323008 251732 323020
rect 251784 323008 251790 323060
rect 277026 322328 277032 322380
rect 277084 322368 277090 322380
rect 407206 322368 407212 322380
rect 277084 322340 407212 322368
rect 277084 322328 277090 322340
rect 407206 322328 407212 322340
rect 407264 322328 407270 322380
rect 291930 322260 291936 322312
rect 291988 322300 291994 322312
rect 483658 322300 483664 322312
rect 291988 322272 483664 322300
rect 291988 322260 291994 322272
rect 483658 322260 483664 322272
rect 483716 322260 483722 322312
rect 288894 322192 288900 322244
rect 288952 322232 288958 322244
rect 528554 322232 528560 322244
rect 288952 322204 528560 322232
rect 288952 322192 288958 322204
rect 528554 322192 528560 322204
rect 528612 322192 528618 322244
rect 283926 321580 283932 321632
rect 283984 321620 283990 321632
rect 284110 321620 284116 321632
rect 283984 321592 284116 321620
rect 283984 321580 283990 321592
rect 284110 321580 284116 321592
rect 284168 321580 284174 321632
rect 3510 320084 3516 320136
rect 3568 320124 3574 320136
rect 234062 320124 234068 320136
rect 3568 320096 234068 320124
rect 3568 320084 3574 320096
rect 234062 320084 234068 320096
rect 234120 320084 234126 320136
rect 252922 319268 252928 319320
rect 252980 319308 252986 319320
rect 253106 319308 253112 319320
rect 252980 319280 253112 319308
rect 252980 319268 252986 319280
rect 253106 319268 253112 319280
rect 253164 319268 253170 319320
rect 316678 313216 316684 313268
rect 316736 313256 316742 313268
rect 580166 313256 580172 313268
rect 316736 313228 580172 313256
rect 316736 313216 316742 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 3510 306280 3516 306332
rect 3568 306320 3574 306332
rect 209038 306320 209044 306332
rect 3568 306292 209044 306320
rect 3568 306280 3574 306292
rect 209038 306280 209044 306292
rect 209096 306280 209102 306332
rect 300210 299412 300216 299464
rect 300268 299452 300274 299464
rect 580166 299452 580172 299464
rect 300268 299424 580172 299452
rect 300268 299412 300274 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 3050 293904 3056 293956
rect 3108 293944 3114 293956
rect 222930 293944 222936 293956
rect 3108 293916 222936 293944
rect 3108 293904 3114 293916
rect 222930 293904 222936 293916
rect 222988 293904 222994 293956
rect 323670 289076 323676 289128
rect 323728 289116 323734 289128
rect 511994 289116 512000 289128
rect 323728 289088 512000 289116
rect 323728 289076 323734 289088
rect 511994 289076 512000 289088
rect 512052 289076 512058 289128
rect 307110 273164 307116 273216
rect 307168 273204 307174 273216
rect 580166 273204 580172 273216
rect 307168 273176 580172 273204
rect 307168 273164 307174 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 3510 267656 3516 267708
rect 3568 267696 3574 267708
rect 232590 267696 232596 267708
rect 3568 267668 232596 267696
rect 3568 267656 3574 267668
rect 232590 267656 232596 267668
rect 232648 267656 232654 267708
rect 314010 259360 314016 259412
rect 314068 259400 314074 259412
rect 580166 259400 580172 259412
rect 314068 259372 580172 259400
rect 314068 259360 314074 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 298830 245556 298836 245608
rect 298888 245596 298894 245608
rect 580166 245596 580172 245608
rect 298888 245568 580172 245596
rect 298888 245556 298894 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 3510 241408 3516 241460
rect 3568 241448 3574 241460
rect 220170 241448 220176 241460
rect 3568 241420 220176 241448
rect 3568 241408 3574 241420
rect 220170 241408 220176 241420
rect 220228 241408 220234 241460
rect 305638 233180 305644 233232
rect 305696 233220 305702 233232
rect 579982 233220 579988 233232
rect 305696 233192 579988 233220
rect 305696 233180 305702 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 231210 215268 231216 215280
rect 3384 215240 231216 215268
rect 3384 215228 3390 215240
rect 231210 215228 231216 215240
rect 231268 215228 231274 215280
rect 295978 206932 295984 206984
rect 296036 206972 296042 206984
rect 579798 206972 579804 206984
rect 296036 206944 579804 206972
rect 296036 206932 296042 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 304258 193128 304264 193180
rect 304316 193168 304322 193180
rect 580166 193168 580172 193180
rect 304316 193140 580172 193168
rect 304316 193128 304322 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 3510 188980 3516 189032
rect 3568 189020 3574 189032
rect 215938 189020 215944 189032
rect 3568 188992 215944 189020
rect 3568 188980 3574 188992
rect 215938 188980 215944 188992
rect 215996 188980 216002 189032
rect 324958 177284 324964 177336
rect 325016 177324 325022 177336
rect 518894 177324 518900 177336
rect 325016 177296 518900 177324
rect 325016 177284 325022 177296
rect 518894 177284 518900 177296
rect 518952 177284 518958 177336
rect 583110 165900 583116 165912
rect 583071 165872 583116 165900
rect 583110 165860 583116 165872
rect 583168 165860 583174 165912
rect 2774 164092 2780 164144
rect 2832 164132 2838 164144
rect 4798 164132 4804 164144
rect 2832 164104 4804 164132
rect 2832 164092 2838 164104
rect 4798 164092 4804 164104
rect 4856 164092 4862 164144
rect 583018 152708 583024 152720
rect 582979 152680 583024 152708
rect 583018 152668 583024 152680
rect 583076 152668 583082 152720
rect 582834 126052 582840 126064
rect 582795 126024 582840 126052
rect 582834 126012 582840 126024
rect 582892 126012 582898 126064
rect 582742 112860 582748 112872
rect 582703 112832 582748 112860
rect 582742 112820 582748 112832
rect 582800 112820 582806 112872
rect 582650 99532 582656 99544
rect 582611 99504 582656 99532
rect 582650 99492 582656 99504
rect 582708 99492 582714 99544
rect 582558 86204 582564 86216
rect 582519 86176 582564 86204
rect 582558 86164 582564 86176
rect 582616 86164 582622 86216
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 214558 85524 214564 85536
rect 3200 85496 214564 85524
rect 3200 85484 3206 85496
rect 214558 85484 214564 85496
rect 214616 85484 214622 85536
rect 582466 73012 582472 73024
rect 582427 72984 582472 73012
rect 582466 72972 582472 72984
rect 582524 72972 582530 73024
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 228450 71720 228456 71732
rect 3476 71692 228456 71720
rect 3476 71680 3482 71692
rect 228450 71680 228456 71692
rect 228508 71680 228514 71732
rect 582374 46356 582380 46368
rect 582335 46328 582380 46356
rect 582374 46316 582380 46328
rect 582432 46316 582438 46368
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 213178 45540 213184 45552
rect 3476 45512 213184 45540
rect 3476 45500 3482 45512
rect 213178 45500 213184 45512
rect 213236 45500 213242 45552
rect 3142 33056 3148 33108
rect 3200 33096 3206 33108
rect 226978 33096 226984 33108
rect 3200 33068 226984 33096
rect 3200 33056 3206 33068
rect 226978 33056 226984 33068
rect 227036 33056 227042 33108
rect 234706 33056 234712 33108
rect 234764 33096 234770 33108
rect 580166 33096 580172 33108
rect 234764 33068 580172 33096
rect 234764 33056 234770 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 294966 20652 294972 20664
rect 3476 20624 294972 20652
rect 3476 20612 3482 20624
rect 294966 20612 294972 20624
rect 295024 20612 295030 20664
rect 157242 17212 157248 17264
rect 157300 17252 157306 17264
rect 250346 17252 250352 17264
rect 157300 17224 250352 17252
rect 157300 17212 157306 17224
rect 250346 17212 250352 17224
rect 250404 17212 250410 17264
rect 327718 17212 327724 17264
rect 327776 17252 327782 17264
rect 550634 17252 550640 17264
rect 327776 17224 550640 17252
rect 327776 17212 327782 17224
rect 550634 17212 550640 17224
rect 550692 17212 550698 17264
rect 267182 15852 267188 15904
rect 267240 15892 267246 15904
rect 316218 15892 316224 15904
rect 267240 15864 316224 15892
rect 267240 15852 267246 15864
rect 316218 15852 316224 15864
rect 316276 15852 316282 15904
rect 323578 15512 323584 15564
rect 323636 15552 323642 15564
rect 327994 15552 328000 15564
rect 323636 15524 328000 15552
rect 323636 15512 323642 15524
rect 327994 15512 328000 15524
rect 328052 15512 328058 15564
rect 215202 14424 215208 14476
rect 215260 14464 215266 14476
rect 222838 14464 222844 14476
rect 215260 14436 222844 14464
rect 215260 14424 215266 14436
rect 222838 14424 222844 14436
rect 222896 14424 222902 14476
rect 287606 13132 287612 13184
rect 287664 13172 287670 13184
rect 517882 13172 517888 13184
rect 287664 13144 517888 13172
rect 287664 13132 287670 13144
rect 517882 13132 517888 13144
rect 517940 13132 517946 13184
rect 5258 13064 5264 13116
rect 5316 13104 5322 13116
rect 173158 13104 173164 13116
rect 5316 13076 173164 13104
rect 5316 13064 5322 13076
rect 173158 13064 173164 13076
rect 173216 13064 173222 13116
rect 228726 13064 228732 13116
rect 228784 13104 228790 13116
rect 233970 13104 233976 13116
rect 228784 13076 233976 13104
rect 228784 13064 228790 13076
rect 233970 13064 233976 13076
rect 234028 13064 234034 13116
rect 292022 13064 292028 13116
rect 292080 13104 292086 13116
rect 556890 13104 556896 13116
rect 292080 13076 556896 13104
rect 292080 13064 292086 13076
rect 556890 13064 556896 13076
rect 556948 13064 556954 13116
rect 280706 12112 280712 12164
rect 280764 12152 280770 12164
rect 442626 12152 442632 12164
rect 280764 12124 442632 12152
rect 280764 12112 280770 12124
rect 442626 12112 442632 12124
rect 442684 12112 442690 12164
rect 280614 12044 280620 12096
rect 280672 12084 280678 12096
rect 445754 12084 445760 12096
rect 280672 12056 445760 12084
rect 280672 12044 280678 12056
rect 445754 12044 445760 12056
rect 445812 12044 445818 12096
rect 280522 11976 280528 12028
rect 280580 12016 280586 12028
rect 448514 12016 448520 12028
rect 280580 11988 448520 12016
rect 280580 11976 280586 11988
rect 448514 11976 448520 11988
rect 448572 11976 448578 12028
rect 281902 11908 281908 11960
rect 281960 11948 281966 11960
rect 453206 11948 453212 11960
rect 281960 11920 453212 11948
rect 281960 11908 281966 11920
rect 453206 11908 453212 11920
rect 453264 11908 453270 11960
rect 281994 11840 282000 11892
rect 282052 11880 282058 11892
rect 456886 11880 456892 11892
rect 282052 11852 456892 11880
rect 282052 11840 282058 11852
rect 456886 11840 456892 11852
rect 456944 11840 456950 11892
rect 165522 11772 165528 11824
rect 165580 11812 165586 11824
rect 224218 11812 224224 11824
rect 165580 11784 224224 11812
rect 165580 11772 165586 11784
rect 224218 11772 224224 11784
rect 224276 11772 224282 11824
rect 282178 11772 282184 11824
rect 282236 11812 282242 11824
rect 459922 11812 459928 11824
rect 282236 11784 459928 11812
rect 282236 11772 282242 11784
rect 459922 11772 459928 11784
rect 459980 11772 459986 11824
rect 65426 11704 65432 11756
rect 65484 11744 65490 11756
rect 240502 11744 240508 11756
rect 65484 11716 240508 11744
rect 65484 11704 65490 11716
rect 240502 11704 240508 11716
rect 240560 11704 240566 11756
rect 282086 11704 282092 11756
rect 282144 11744 282150 11756
rect 463970 11744 463976 11756
rect 282144 11716 463976 11744
rect 282144 11704 282150 11716
rect 463970 11704 463976 11716
rect 464028 11704 464034 11756
rect 324406 11636 324412 11688
rect 324464 11676 324470 11688
rect 325602 11676 325608 11688
rect 324464 11648 325608 11676
rect 324464 11636 324470 11648
rect 325602 11636 325608 11648
rect 325660 11636 325666 11688
rect 407206 11636 407212 11688
rect 407264 11676 407270 11688
rect 408402 11676 408408 11688
rect 407264 11648 408408 11676
rect 407264 11636 407270 11648
rect 408402 11636 408408 11648
rect 408460 11636 408466 11688
rect 423766 11636 423772 11688
rect 423824 11676 423830 11688
rect 424962 11676 424968 11688
rect 423824 11648 424968 11676
rect 423824 11636 423830 11648
rect 424962 11636 424968 11648
rect 425020 11636 425026 11688
rect 272702 10956 272708 11008
rect 272760 10996 272766 11008
rect 367738 10996 367744 11008
rect 272760 10968 367744 10996
rect 272760 10956 272766 10968
rect 367738 10956 367744 10968
rect 367796 10956 367802 11008
rect 272610 10888 272616 10940
rect 272668 10928 272674 10940
rect 371234 10928 371240 10940
rect 272668 10900 371240 10928
rect 272668 10888 272674 10900
rect 371234 10888 371240 10900
rect 371292 10888 371298 10940
rect 273990 10820 273996 10872
rect 274048 10860 274054 10872
rect 373994 10860 374000 10872
rect 274048 10832 374000 10860
rect 274048 10820 274054 10832
rect 373994 10820 374000 10832
rect 374052 10820 374058 10872
rect 274174 10752 274180 10804
rect 274232 10792 274238 10804
rect 378410 10792 378416 10804
rect 274232 10764 378416 10792
rect 274232 10752 274238 10764
rect 378410 10752 378416 10764
rect 378468 10752 378474 10804
rect 274082 10684 274088 10736
rect 274140 10724 274146 10736
rect 382366 10724 382372 10736
rect 274140 10696 382372 10724
rect 274140 10684 274146 10696
rect 382366 10684 382372 10696
rect 382424 10684 382430 10736
rect 275462 10616 275468 10668
rect 275520 10656 275526 10668
rect 385586 10656 385592 10668
rect 275520 10628 385592 10656
rect 275520 10616 275526 10628
rect 385586 10616 385592 10628
rect 385644 10616 385650 10668
rect 275370 10548 275376 10600
rect 275428 10588 275434 10600
rect 389450 10588 389456 10600
rect 275428 10560 389456 10588
rect 275428 10548 275434 10560
rect 389450 10548 389456 10560
rect 389508 10548 389514 10600
rect 150342 10480 150348 10532
rect 150400 10520 150406 10532
rect 250162 10520 250168 10532
rect 150400 10492 250168 10520
rect 150400 10480 150406 10492
rect 250162 10480 250168 10492
rect 250220 10480 250226 10532
rect 275646 10480 275652 10532
rect 275704 10520 275710 10532
rect 392578 10520 392584 10532
rect 275704 10492 392584 10520
rect 275704 10480 275710 10492
rect 392578 10480 392584 10492
rect 392636 10480 392642 10532
rect 122742 10412 122748 10464
rect 122800 10452 122806 10464
rect 247494 10452 247500 10464
rect 122800 10424 247500 10452
rect 122800 10412 122806 10424
rect 247494 10412 247500 10424
rect 247552 10412 247558 10464
rect 275278 10412 275284 10464
rect 275336 10452 275342 10464
rect 396074 10452 396080 10464
rect 275336 10424 396080 10452
rect 275336 10412 275342 10424
rect 396074 10412 396080 10424
rect 396132 10412 396138 10464
rect 119798 10344 119804 10396
rect 119856 10384 119862 10396
rect 247402 10384 247408 10396
rect 119856 10356 247408 10384
rect 119856 10344 119862 10356
rect 247402 10344 247408 10356
rect 247460 10344 247466 10396
rect 276566 10344 276572 10396
rect 276624 10384 276630 10396
rect 400122 10384 400128 10396
rect 276624 10356 400128 10384
rect 276624 10344 276630 10356
rect 400122 10344 400128 10356
rect 400180 10344 400186 10396
rect 115842 10276 115848 10328
rect 115900 10316 115906 10328
rect 246390 10316 246396 10328
rect 115900 10288 246396 10316
rect 115900 10276 115906 10288
rect 246390 10276 246396 10288
rect 246448 10276 246454 10328
rect 277118 10276 277124 10328
rect 277176 10316 277182 10328
rect 403526 10316 403532 10328
rect 277176 10288 403532 10316
rect 277176 10276 277182 10288
rect 403526 10276 403532 10288
rect 403584 10276 403590 10328
rect 272518 10208 272524 10260
rect 272576 10248 272582 10260
rect 364610 10248 364616 10260
rect 272576 10220 364616 10248
rect 272576 10208 272582 10220
rect 364610 10208 364616 10220
rect 364668 10208 364674 10260
rect 272794 10140 272800 10192
rect 272852 10180 272858 10192
rect 360746 10180 360752 10192
rect 272852 10152 360752 10180
rect 272852 10140 272858 10152
rect 360746 10140 360752 10152
rect 360804 10140 360810 10192
rect 271138 10072 271144 10124
rect 271196 10112 271202 10124
rect 357526 10112 357532 10124
rect 271196 10084 357532 10112
rect 271196 10072 271202 10084
rect 357526 10072 357532 10084
rect 357584 10072 357590 10124
rect 271414 10004 271420 10056
rect 271472 10044 271478 10056
rect 353570 10044 353576 10056
rect 271472 10016 353576 10044
rect 271472 10004 271478 10016
rect 353570 10004 353576 10016
rect 353628 10004 353634 10056
rect 270586 9936 270592 9988
rect 270644 9976 270650 9988
rect 350442 9976 350448 9988
rect 270644 9948 350448 9976
rect 270644 9936 270650 9948
rect 350442 9936 350448 9948
rect 350500 9936 350506 9988
rect 271322 9868 271328 9920
rect 271380 9908 271386 9920
rect 346946 9908 346952 9920
rect 271380 9880 346952 9908
rect 271380 9868 271386 9880
rect 346946 9868 346952 9880
rect 347004 9868 347010 9920
rect 270034 9800 270040 9852
rect 270092 9840 270098 9852
rect 342898 9840 342904 9852
rect 270092 9812 342904 9840
rect 270092 9800 270098 9812
rect 342898 9800 342904 9812
rect 342956 9800 342962 9852
rect 270126 9732 270132 9784
rect 270184 9772 270190 9784
rect 339494 9772 339500 9784
rect 270184 9744 339500 9772
rect 270184 9732 270190 9744
rect 339494 9732 339500 9744
rect 339552 9732 339558 9784
rect 231026 9392 231032 9444
rect 231084 9432 231090 9444
rect 257430 9432 257436 9444
rect 231084 9404 257436 9432
rect 231084 9392 231090 9404
rect 257430 9392 257436 9404
rect 257488 9392 257494 9444
rect 160094 9324 160100 9376
rect 160152 9364 160158 9376
rect 251542 9364 251548 9376
rect 160152 9336 251548 9364
rect 160152 9324 160158 9336
rect 251542 9324 251548 9336
rect 251600 9324 251606 9376
rect 266078 9324 266084 9376
rect 266136 9364 266142 9376
rect 297266 9364 297272 9376
rect 266136 9336 297272 9364
rect 266136 9324 266142 9336
rect 297266 9324 297272 9336
rect 297324 9324 297330 9376
rect 142430 9256 142436 9308
rect 142488 9296 142494 9308
rect 249242 9296 249248 9308
rect 142488 9268 249248 9296
rect 142488 9256 142494 9268
rect 249242 9256 249248 9268
rect 249300 9256 249306 9308
rect 265986 9256 265992 9308
rect 266044 9296 266050 9308
rect 300762 9296 300768 9308
rect 266044 9268 300768 9296
rect 266044 9256 266050 9268
rect 300762 9256 300768 9268
rect 300820 9256 300826 9308
rect 138842 9188 138848 9240
rect 138900 9228 138906 9240
rect 248690 9228 248696 9240
rect 138900 9200 248696 9228
rect 138900 9188 138906 9200
rect 248690 9188 248696 9200
rect 248748 9188 248754 9240
rect 265894 9188 265900 9240
rect 265952 9228 265958 9240
rect 304350 9228 304356 9240
rect 265952 9200 304356 9228
rect 265952 9188 265958 9200
rect 304350 9188 304356 9200
rect 304408 9188 304414 9240
rect 135254 9120 135260 9172
rect 135312 9160 135318 9172
rect 248966 9160 248972 9172
rect 135312 9132 248972 9160
rect 135312 9120 135318 9132
rect 248966 9120 248972 9132
rect 249024 9120 249030 9172
rect 268470 9120 268476 9172
rect 268528 9160 268534 9172
rect 326798 9160 326804 9172
rect 268528 9132 326804 9160
rect 268528 9120 268534 9132
rect 326798 9120 326804 9132
rect 326856 9120 326862 9172
rect 83274 9052 83280 9104
rect 83332 9092 83338 9104
rect 243354 9092 243360 9104
rect 83332 9064 243360 9092
rect 83332 9052 83338 9064
rect 243354 9052 243360 9064
rect 243412 9052 243418 9104
rect 284478 9052 284484 9104
rect 284536 9092 284542 9104
rect 489914 9092 489920 9104
rect 284536 9064 489920 9092
rect 284536 9052 284542 9064
rect 489914 9052 489920 9064
rect 489972 9052 489978 9104
rect 79686 8984 79692 9036
rect 79744 9024 79750 9036
rect 243262 9024 243268 9036
rect 79744 8996 243268 9024
rect 79744 8984 79750 8996
rect 243262 8984 243268 8996
rect 243320 8984 243326 9036
rect 294782 8984 294788 9036
rect 294840 9024 294846 9036
rect 573910 9024 573916 9036
rect 294840 8996 573916 9024
rect 294840 8984 294846 8996
rect 573910 8984 573916 8996
rect 573968 8984 573974 9036
rect 8754 8916 8760 8968
rect 8812 8956 8818 8968
rect 235350 8956 235356 8968
rect 8812 8928 235356 8956
rect 8812 8916 8818 8928
rect 235350 8916 235356 8928
rect 235408 8916 235414 8968
rect 294690 8916 294696 8968
rect 294748 8956 294754 8968
rect 577406 8956 577412 8968
rect 294748 8928 577412 8956
rect 294748 8916 294754 8928
rect 577406 8916 577412 8928
rect 577464 8916 577470 8968
rect 199102 8168 199108 8220
rect 199160 8208 199166 8220
rect 255958 8208 255964 8220
rect 199160 8180 255964 8208
rect 199160 8168 199166 8180
rect 255958 8168 255964 8180
rect 256016 8168 256022 8220
rect 181438 8100 181444 8152
rect 181496 8140 181502 8152
rect 252922 8140 252928 8152
rect 181496 8112 252928 8140
rect 181496 8100 181502 8112
rect 252922 8100 252928 8112
rect 252980 8100 252986 8152
rect 174262 8032 174268 8084
rect 174320 8072 174326 8084
rect 253014 8072 253020 8084
rect 174320 8044 253020 8072
rect 174320 8032 174326 8044
rect 253014 8032 253020 8044
rect 253072 8032 253078 8084
rect 170766 7964 170772 8016
rect 170824 8004 170830 8016
rect 251634 8004 251640 8016
rect 170824 7976 251640 8004
rect 170824 7964 170830 7976
rect 251634 7964 251640 7976
rect 251692 7964 251698 8016
rect 280982 7964 280988 8016
rect 281040 8004 281046 8016
rect 441522 8004 441528 8016
rect 281040 7976 441528 8004
rect 281040 7964 281046 7976
rect 441522 7964 441528 7976
rect 441580 7964 441586 8016
rect 167178 7896 167184 7948
rect 167236 7936 167242 7948
rect 252002 7936 252008 7948
rect 167236 7908 252008 7936
rect 167236 7896 167242 7908
rect 252002 7896 252008 7908
rect 252060 7896 252066 7948
rect 280890 7896 280896 7948
rect 280948 7936 280954 7948
rect 445018 7936 445024 7948
rect 280948 7908 445024 7936
rect 280948 7896 280954 7908
rect 445018 7896 445024 7908
rect 445076 7896 445082 7948
rect 163682 7828 163688 7880
rect 163740 7868 163746 7880
rect 251358 7868 251364 7880
rect 163740 7840 251364 7868
rect 163740 7828 163746 7840
rect 251358 7828 251364 7840
rect 251416 7828 251422 7880
rect 281074 7828 281080 7880
rect 281132 7868 281138 7880
rect 448606 7868 448612 7880
rect 281132 7840 448612 7868
rect 281132 7828 281138 7840
rect 448606 7828 448612 7840
rect 448664 7828 448670 7880
rect 158898 7760 158904 7812
rect 158956 7800 158962 7812
rect 251450 7800 251456 7812
rect 158956 7772 251456 7800
rect 158956 7760 158962 7772
rect 251450 7760 251456 7772
rect 251508 7760 251514 7812
rect 280798 7760 280804 7812
rect 280856 7800 280862 7812
rect 452102 7800 452108 7812
rect 280856 7772 452108 7800
rect 280856 7760 280862 7772
rect 452102 7760 452108 7772
rect 452160 7760 452166 7812
rect 131758 7692 131764 7744
rect 131816 7732 131822 7744
rect 248782 7732 248788 7744
rect 131816 7704 248788 7732
rect 131816 7692 131822 7704
rect 248782 7692 248788 7704
rect 248840 7692 248846 7744
rect 282270 7692 282276 7744
rect 282328 7732 282334 7744
rect 455690 7732 455696 7744
rect 282328 7704 455696 7732
rect 282328 7692 282334 7704
rect 455690 7692 455696 7704
rect 455748 7692 455754 7744
rect 128170 7624 128176 7676
rect 128228 7664 128234 7676
rect 247310 7664 247316 7676
rect 128228 7636 247316 7664
rect 128228 7624 128234 7636
rect 247310 7624 247316 7636
rect 247368 7624 247374 7676
rect 282454 7624 282460 7676
rect 282512 7664 282518 7676
rect 459186 7664 459192 7676
rect 282512 7636 459192 7664
rect 282512 7624 282518 7636
rect 459186 7624 459192 7636
rect 459244 7624 459250 7676
rect 9950 7556 9956 7608
rect 10008 7596 10014 7608
rect 177298 7596 177304 7608
rect 10008 7568 177304 7596
rect 10008 7556 10014 7568
rect 177298 7556 177304 7568
rect 177356 7556 177362 7608
rect 177850 7556 177856 7608
rect 177908 7596 177914 7608
rect 253106 7596 253112 7608
rect 177908 7568 253112 7596
rect 177908 7556 177914 7568
rect 253106 7556 253112 7568
rect 253164 7556 253170 7608
rect 282362 7556 282368 7608
rect 282420 7596 282426 7608
rect 462774 7596 462780 7608
rect 282420 7568 462780 7596
rect 282420 7556 282426 7568
rect 462774 7556 462780 7568
rect 462832 7556 462838 7608
rect 234614 6808 234620 6860
rect 234672 6848 234678 6860
rect 580166 6848 580172 6860
rect 234672 6820 580172 6848
rect 234672 6808 234678 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 3326 6740 3332 6792
rect 3384 6780 3390 6792
rect 294598 6780 294604 6792
rect 3384 6752 294604 6780
rect 3384 6740 3390 6752
rect 294598 6740 294604 6752
rect 294656 6740 294662 6792
rect 208578 6672 208584 6724
rect 208636 6712 208642 6724
rect 255866 6712 255872 6724
rect 208636 6684 255872 6712
rect 208636 6672 208642 6684
rect 255866 6672 255872 6684
rect 255924 6672 255930 6724
rect 271598 6672 271604 6724
rect 271656 6712 271662 6724
rect 356330 6712 356336 6724
rect 271656 6684 356336 6712
rect 271656 6672 271662 6684
rect 356330 6672 356336 6684
rect 356388 6672 356394 6724
rect 205082 6604 205088 6656
rect 205140 6644 205146 6656
rect 255682 6644 255688 6656
rect 205140 6616 255688 6644
rect 205140 6604 205146 6616
rect 255682 6604 255688 6616
rect 255740 6604 255746 6656
rect 273070 6604 273076 6656
rect 273128 6644 273134 6656
rect 359918 6644 359924 6656
rect 273128 6616 359924 6644
rect 273128 6604 273134 6616
rect 359918 6604 359924 6616
rect 359976 6604 359982 6656
rect 201494 6536 201500 6588
rect 201552 6576 201558 6588
rect 255774 6576 255780 6588
rect 201552 6548 255780 6576
rect 201552 6536 201558 6548
rect 255774 6536 255780 6548
rect 255832 6536 255838 6588
rect 272978 6536 272984 6588
rect 273036 6576 273042 6588
rect 363506 6576 363512 6588
rect 273036 6548 363512 6576
rect 273036 6536 273042 6548
rect 363506 6536 363512 6548
rect 363564 6536 363570 6588
rect 183738 6468 183744 6520
rect 183796 6508 183802 6520
rect 252830 6508 252836 6520
rect 183796 6480 252836 6508
rect 183796 6468 183802 6480
rect 252830 6468 252836 6480
rect 252888 6468 252894 6520
rect 273162 6468 273168 6520
rect 273220 6508 273226 6520
rect 367002 6508 367008 6520
rect 273220 6480 367008 6508
rect 273220 6468 273226 6480
rect 367002 6468 367008 6480
rect 367060 6468 367066 6520
rect 176654 6400 176660 6452
rect 176712 6440 176718 6452
rect 253382 6440 253388 6452
rect 176712 6412 253388 6440
rect 176712 6400 176718 6412
rect 253382 6400 253388 6412
rect 253440 6400 253446 6452
rect 272886 6400 272892 6452
rect 272944 6440 272950 6452
rect 370590 6440 370596 6452
rect 272944 6412 370596 6440
rect 272944 6400 272950 6412
rect 370590 6400 370596 6412
rect 370648 6400 370654 6452
rect 102226 6332 102232 6384
rect 102284 6372 102290 6384
rect 180058 6372 180064 6384
rect 102284 6344 180064 6372
rect 102284 6332 102290 6344
rect 180058 6332 180064 6344
rect 180116 6332 180122 6384
rect 180242 6332 180248 6384
rect 180300 6372 180306 6384
rect 253658 6372 253664 6384
rect 180300 6344 253664 6372
rect 180300 6332 180306 6344
rect 253658 6332 253664 6344
rect 253716 6332 253722 6384
rect 274266 6332 274272 6384
rect 274324 6372 274330 6384
rect 374086 6372 374092 6384
rect 274324 6344 374092 6372
rect 274324 6332 274330 6344
rect 374086 6332 374092 6344
rect 374144 6332 374150 6384
rect 173158 6264 173164 6316
rect 173216 6304 173222 6316
rect 252738 6304 252744 6316
rect 173216 6276 252744 6304
rect 173216 6264 173222 6276
rect 252738 6264 252744 6276
rect 252796 6264 252802 6316
rect 273714 6264 273720 6316
rect 273772 6304 273778 6316
rect 377674 6304 377680 6316
rect 273772 6276 377680 6304
rect 273772 6264 273778 6276
rect 377674 6264 377680 6276
rect 377732 6264 377738 6316
rect 28810 6196 28816 6248
rect 28868 6236 28874 6248
rect 130378 6236 130384 6248
rect 28868 6208 130384 6236
rect 28868 6196 28874 6208
rect 130378 6196 130384 6208
rect 130436 6196 130442 6248
rect 130562 6196 130568 6248
rect 130620 6236 130626 6248
rect 247218 6236 247224 6248
rect 130620 6208 247224 6236
rect 130620 6196 130626 6208
rect 247218 6196 247224 6208
rect 247276 6196 247282 6248
rect 273898 6196 273904 6248
rect 273956 6236 273962 6248
rect 381170 6236 381176 6248
rect 273956 6208 381176 6236
rect 273956 6196 273962 6208
rect 381170 6196 381176 6208
rect 381228 6196 381234 6248
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 235258 6168 235264 6180
rect 4120 6140 235264 6168
rect 4120 6128 4126 6140
rect 235258 6128 235264 6140
rect 235316 6128 235322 6180
rect 266998 6128 267004 6180
rect 267056 6168 267062 6180
rect 273622 6168 273628 6180
rect 267056 6140 273628 6168
rect 267056 6128 267062 6140
rect 273622 6128 273628 6140
rect 273680 6128 273686 6180
rect 273806 6128 273812 6180
rect 273864 6168 273870 6180
rect 384758 6168 384764 6180
rect 273864 6140 384764 6168
rect 273864 6128 273870 6140
rect 384758 6128 384764 6140
rect 384816 6128 384822 6180
rect 271506 6060 271512 6112
rect 271564 6100 271570 6112
rect 352834 6100 352840 6112
rect 271564 6072 352840 6100
rect 271564 6060 271570 6072
rect 352834 6060 352840 6072
rect 352892 6060 352898 6112
rect 271046 5992 271052 6044
rect 271104 6032 271110 6044
rect 349246 6032 349252 6044
rect 271104 6004 349252 6032
rect 271104 5992 271110 6004
rect 349246 5992 349252 6004
rect 349304 5992 349310 6044
rect 270954 5924 270960 5976
rect 271012 5964 271018 5976
rect 345750 5964 345756 5976
rect 271012 5936 345756 5964
rect 271012 5924 271018 5936
rect 345750 5924 345756 5936
rect 345808 5924 345814 5976
rect 269850 5856 269856 5908
rect 269908 5896 269914 5908
rect 342162 5896 342168 5908
rect 269908 5868 342168 5896
rect 269908 5856 269914 5868
rect 342162 5856 342168 5868
rect 342220 5856 342226 5908
rect 269942 5788 269948 5840
rect 270000 5828 270006 5840
rect 338666 5828 338672 5840
rect 270000 5800 338672 5828
rect 270000 5788 270006 5800
rect 338666 5788 338672 5800
rect 338724 5788 338730 5840
rect 269666 5720 269672 5772
rect 269724 5760 269730 5772
rect 335078 5760 335084 5772
rect 269724 5732 335084 5760
rect 269724 5720 269730 5732
rect 335078 5720 335084 5732
rect 335136 5720 335142 5772
rect 268654 5652 268660 5704
rect 268712 5692 268718 5704
rect 331582 5692 331588 5704
rect 268712 5664 331588 5692
rect 268712 5652 268718 5664
rect 331582 5652 331588 5664
rect 331640 5652 331646 5704
rect 196802 5516 196808 5568
rect 196860 5556 196866 5568
rect 202138 5556 202144 5568
rect 196860 5528 202144 5556
rect 196860 5516 196866 5528
rect 202138 5516 202144 5528
rect 202196 5516 202202 5568
rect 218054 5448 218060 5500
rect 218112 5488 218118 5500
rect 232498 5488 232504 5500
rect 218112 5460 232504 5488
rect 218112 5448 218118 5460
rect 232498 5448 232504 5460
rect 232556 5448 232562 5500
rect 233050 5448 233056 5500
rect 233108 5488 233114 5500
rect 253474 5488 253480 5500
rect 233108 5460 253480 5488
rect 233108 5448 233114 5460
rect 253474 5448 253480 5460
rect 253532 5448 253538 5500
rect 253842 5448 253848 5500
rect 253900 5488 253906 5500
rect 267734 5488 267740 5500
rect 253900 5460 267740 5488
rect 253900 5448 253906 5460
rect 267734 5448 267740 5460
rect 267792 5448 267798 5500
rect 272426 5448 272432 5500
rect 272484 5488 272490 5500
rect 284386 5488 284392 5500
rect 272484 5460 284392 5488
rect 272484 5448 272490 5460
rect 284386 5448 284392 5460
rect 284444 5448 284450 5500
rect 288986 5448 288992 5500
rect 289044 5488 289050 5500
rect 289538 5488 289544 5500
rect 289044 5460 289544 5488
rect 289044 5448 289050 5460
rect 289538 5448 289544 5460
rect 289596 5448 289602 5500
rect 189718 5380 189724 5432
rect 189776 5420 189782 5432
rect 233878 5420 233884 5432
rect 189776 5392 233884 5420
rect 189776 5380 189782 5392
rect 233878 5380 233884 5392
rect 233936 5380 233942 5432
rect 240502 5380 240508 5432
rect 240560 5420 240566 5432
rect 258718 5420 258724 5432
rect 240560 5392 258724 5420
rect 240560 5380 240566 5392
rect 258718 5380 258724 5392
rect 258776 5380 258782 5432
rect 263134 5380 263140 5432
rect 263192 5420 263198 5432
rect 276014 5420 276020 5432
rect 263192 5392 276020 5420
rect 263192 5380 263198 5392
rect 276014 5380 276020 5392
rect 276072 5380 276078 5432
rect 186130 5312 186136 5364
rect 186188 5352 186194 5364
rect 204898 5352 204904 5364
rect 186188 5324 204904 5352
rect 186188 5312 186194 5324
rect 204898 5312 204904 5324
rect 204956 5312 204962 5364
rect 211062 5312 211068 5364
rect 211120 5352 211126 5364
rect 255406 5352 255412 5364
rect 211120 5324 255412 5352
rect 211120 5312 211126 5324
rect 255406 5312 255412 5324
rect 255464 5312 255470 5364
rect 262490 5312 262496 5364
rect 262548 5352 262554 5364
rect 278314 5352 278320 5364
rect 262548 5324 278320 5352
rect 262548 5312 262554 5324
rect 278314 5312 278320 5324
rect 278372 5312 278378 5364
rect 171962 5244 171968 5296
rect 172020 5284 172026 5296
rect 206278 5284 206284 5296
rect 172020 5256 206284 5284
rect 172020 5244 172026 5256
rect 206278 5244 206284 5256
rect 206336 5244 206342 5296
rect 207382 5244 207388 5296
rect 207440 5284 207446 5296
rect 255590 5284 255596 5296
rect 207440 5256 255596 5284
rect 207440 5244 207446 5256
rect 255590 5244 255596 5256
rect 255648 5244 255654 5296
rect 264422 5244 264428 5296
rect 264480 5284 264486 5296
rect 279510 5284 279516 5296
rect 264480 5256 279516 5284
rect 264480 5244 264486 5256
rect 279510 5244 279516 5256
rect 279568 5244 279574 5296
rect 182542 5176 182548 5228
rect 182600 5216 182606 5228
rect 196618 5216 196624 5228
rect 182600 5188 196624 5216
rect 182600 5176 182606 5188
rect 196618 5176 196624 5188
rect 196676 5176 196682 5228
rect 203886 5176 203892 5228
rect 203944 5216 203950 5228
rect 256050 5216 256056 5228
rect 203944 5188 256056 5216
rect 203944 5176 203950 5188
rect 256050 5176 256056 5188
rect 256108 5176 256114 5228
rect 264514 5176 264520 5228
rect 264572 5216 264578 5228
rect 281902 5216 281908 5228
rect 264572 5188 281908 5216
rect 264572 5176 264578 5188
rect 281902 5176 281908 5188
rect 281960 5176 281966 5228
rect 376110 5176 376116 5228
rect 376168 5216 376174 5228
rect 402514 5216 402520 5228
rect 376168 5188 402520 5216
rect 376168 5176 376174 5188
rect 402514 5176 402520 5188
rect 402572 5176 402578 5228
rect 175458 5108 175464 5160
rect 175516 5148 175522 5160
rect 197998 5148 198004 5160
rect 175516 5120 198004 5148
rect 175516 5108 175522 5120
rect 197998 5108 198004 5120
rect 198056 5108 198062 5160
rect 200298 5108 200304 5160
rect 200356 5148 200362 5160
rect 255498 5148 255504 5160
rect 200356 5120 255504 5148
rect 200356 5108 200362 5120
rect 255498 5108 255504 5120
rect 255556 5108 255562 5160
rect 264330 5108 264336 5160
rect 264388 5148 264394 5160
rect 283098 5148 283104 5160
rect 264388 5120 283104 5148
rect 264388 5108 264394 5120
rect 283098 5108 283104 5120
rect 283156 5108 283162 5160
rect 335998 5108 336004 5160
rect 336056 5148 336062 5160
rect 391842 5148 391848 5160
rect 336056 5120 391848 5148
rect 336056 5108 336062 5120
rect 391842 5108 391848 5120
rect 391900 5108 391906 5160
rect 393958 5108 393964 5160
rect 394016 5148 394022 5160
rect 409598 5148 409604 5160
rect 394016 5120 409604 5148
rect 394016 5108 394022 5120
rect 409598 5108 409604 5120
rect 409656 5108 409662 5160
rect 129366 5040 129372 5092
rect 129424 5080 129430 5092
rect 247126 5080 247132 5092
rect 129424 5052 247132 5080
rect 129424 5040 129430 5052
rect 247126 5040 247132 5052
rect 247184 5040 247190 5092
rect 264606 5040 264612 5092
rect 264664 5080 264670 5092
rect 285398 5080 285404 5092
rect 264664 5052 285404 5080
rect 264664 5040 264670 5052
rect 285398 5040 285404 5052
rect 285456 5040 285462 5092
rect 286318 5040 286324 5092
rect 286376 5080 286382 5092
rect 309042 5080 309048 5092
rect 286376 5052 309048 5080
rect 286376 5040 286382 5052
rect 309042 5040 309048 5052
rect 309100 5040 309106 5092
rect 331858 5040 331864 5092
rect 331916 5080 331922 5092
rect 495894 5080 495900 5092
rect 331916 5052 495900 5080
rect 331916 5040 331922 5052
rect 495894 5040 495900 5052
rect 495952 5040 495958 5092
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 7708 4984 232176 5012
rect 7708 4972 7714 4984
rect 2866 4904 2872 4956
rect 2924 4944 2930 4956
rect 232041 4947 232099 4953
rect 232041 4944 232053 4947
rect 2924 4916 232053 4944
rect 2924 4904 2930 4916
rect 232041 4913 232053 4916
rect 232087 4913 232099 4947
rect 232148 4944 232176 4984
rect 234614 4972 234620 5024
rect 234672 5012 234678 5024
rect 254578 5012 254584 5024
rect 234672 4984 254584 5012
rect 234672 4972 234678 4984
rect 254578 4972 254584 4984
rect 254636 4972 254642 5024
rect 264698 4972 264704 5024
rect 264756 5012 264762 5024
rect 286594 5012 286600 5024
rect 264756 4984 286600 5012
rect 264756 4972 264762 4984
rect 286594 4972 286600 4984
rect 286652 4972 286658 5024
rect 298738 4972 298744 5024
rect 298796 5012 298802 5024
rect 298796 4984 320772 5012
rect 298796 4972 298802 4984
rect 235166 4944 235172 4956
rect 232148 4916 235172 4944
rect 232041 4907 232099 4913
rect 235166 4904 235172 4916
rect 235224 4904 235230 4956
rect 238110 4904 238116 4956
rect 238168 4944 238174 4956
rect 258350 4944 258356 4956
rect 238168 4916 258356 4944
rect 238168 4904 238174 4916
rect 258350 4904 258356 4916
rect 258408 4904 258414 4956
rect 267274 4904 267280 4956
rect 267332 4944 267338 4956
rect 319714 4944 319720 4956
rect 267332 4916 319720 4944
rect 267332 4904 267338 4916
rect 319714 4904 319720 4916
rect 319772 4904 319778 4956
rect 320744 4944 320772 4984
rect 320818 4972 320824 5024
rect 320876 5012 320882 5024
rect 494698 5012 494704 5024
rect 320876 4984 494704 5012
rect 320876 4972 320882 4984
rect 494698 4972 494704 4984
rect 494756 4972 494762 5024
rect 320910 4944 320916 4956
rect 320744 4916 320916 4944
rect 320910 4904 320916 4916
rect 320968 4904 320974 4956
rect 322198 4904 322204 4956
rect 322256 4944 322262 4956
rect 505370 4944 505376 4956
rect 322256 4916 505376 4944
rect 322256 4904 322262 4916
rect 505370 4904 505376 4916
rect 505428 4904 505434 4956
rect 1670 4836 1676 4888
rect 1728 4876 1734 4888
rect 234890 4876 234896 4888
rect 1728 4848 234896 4876
rect 1728 4836 1734 4848
rect 234890 4836 234896 4848
rect 234948 4836 234954 4888
rect 239306 4836 239312 4888
rect 239364 4876 239370 4888
rect 259730 4876 259736 4888
rect 239364 4848 259736 4876
rect 239364 4836 239370 4848
rect 259730 4836 259736 4848
rect 259788 4836 259794 4888
rect 264146 4836 264152 4888
rect 264204 4876 264210 4888
rect 288986 4876 288992 4888
rect 264204 4848 288992 4876
rect 264204 4836 264210 4848
rect 288986 4836 288992 4848
rect 289044 4836 289050 4888
rect 289538 4836 289544 4888
rect 289596 4876 289602 4888
rect 532510 4876 532516 4888
rect 289596 4848 532516 4876
rect 289596 4836 289602 4848
rect 532510 4836 532516 4848
rect 532568 4836 532574 4888
rect 566 4768 572 4820
rect 624 4808 630 4820
rect 232041 4811 232099 4817
rect 624 4780 231992 4808
rect 624 4768 630 4780
rect 221550 4700 221556 4752
rect 221608 4740 221614 4752
rect 231118 4740 231124 4752
rect 221608 4712 231124 4740
rect 221608 4700 221614 4712
rect 231118 4700 231124 4712
rect 231176 4700 231182 4752
rect 231964 4740 231992 4780
rect 232041 4777 232053 4811
rect 232087 4808 232099 4811
rect 235074 4808 235080 4820
rect 232087 4780 235080 4808
rect 232087 4777 232099 4780
rect 232041 4771 232099 4777
rect 235074 4768 235080 4780
rect 235132 4768 235138 4820
rect 237006 4768 237012 4820
rect 237064 4808 237070 4820
rect 258626 4808 258632 4820
rect 237064 4780 258632 4808
rect 237064 4768 237070 4780
rect 258626 4768 258632 4780
rect 258684 4768 258690 4820
rect 265802 4768 265808 4820
rect 265860 4808 265866 4820
rect 292574 4808 292580 4820
rect 265860 4780 292580 4808
rect 265860 4768 265866 4780
rect 292574 4768 292580 4780
rect 292632 4768 292638 4820
rect 294966 4768 294972 4820
rect 295024 4808 295030 4820
rect 576302 4808 576308 4820
rect 295024 4780 576308 4808
rect 295024 4768 295030 4780
rect 576302 4768 576308 4780
rect 576360 4768 576366 4820
rect 234982 4740 234988 4752
rect 231964 4712 234988 4740
rect 234982 4700 234988 4712
rect 235040 4700 235046 4752
rect 249978 4740 249984 4752
rect 238726 4712 249984 4740
rect 231670 4632 231676 4684
rect 231728 4672 231734 4684
rect 238726 4672 238754 4712
rect 249978 4700 249984 4712
rect 250036 4700 250042 4752
rect 263042 4700 263048 4752
rect 263100 4740 263106 4752
rect 274818 4740 274824 4752
rect 263100 4712 274824 4740
rect 263100 4700 263106 4712
rect 274818 4700 274824 4712
rect 274876 4700 274882 4752
rect 231728 4644 238754 4672
rect 231728 4632 231734 4644
rect 241698 4632 241704 4684
rect 241756 4672 241762 4684
rect 258810 4672 258816 4684
rect 241756 4644 258816 4672
rect 241756 4632 241762 4644
rect 258810 4632 258816 4644
rect 258868 4632 258874 4684
rect 262950 4632 262956 4684
rect 263008 4672 263014 4684
rect 271230 4672 271236 4684
rect 263008 4644 271236 4672
rect 263008 4632 263014 4644
rect 271230 4632 271236 4644
rect 271288 4632 271294 4684
rect 242894 4564 242900 4616
rect 242952 4604 242958 4616
rect 259822 4604 259828 4616
rect 242952 4576 259828 4604
rect 242952 4564 242958 4576
rect 259822 4564 259828 4576
rect 259880 4564 259886 4616
rect 231762 4496 231768 4548
rect 231820 4536 231826 4548
rect 247586 4536 247592 4548
rect 231820 4508 247592 4536
rect 231820 4496 231826 4508
rect 247586 4496 247592 4508
rect 247644 4496 247650 4548
rect 246390 4428 246396 4480
rect 246448 4468 246454 4480
rect 259638 4468 259644 4480
rect 246448 4440 259644 4468
rect 246448 4428 246454 4440
rect 259638 4428 259644 4440
rect 259696 4428 259702 4480
rect 244090 4360 244096 4412
rect 244148 4400 244154 4412
rect 251818 4400 251824 4412
rect 244148 4372 251824 4400
rect 244148 4360 244154 4372
rect 251818 4360 251824 4372
rect 251876 4360 251882 4412
rect 277118 4360 277124 4412
rect 277176 4400 277182 4412
rect 277670 4400 277676 4412
rect 277176 4372 277676 4400
rect 277176 4360 277182 4372
rect 277670 4360 277676 4372
rect 277728 4360 277734 4412
rect 290182 4292 290188 4344
rect 290240 4332 290246 4344
rect 295426 4332 295432 4344
rect 290240 4304 295432 4332
rect 290240 4292 290246 4304
rect 295426 4292 295432 4304
rect 295484 4292 295490 4344
rect 293678 4224 293684 4276
rect 293736 4264 293742 4276
rect 295518 4264 295524 4276
rect 293736 4236 295524 4264
rect 293736 4224 293742 4236
rect 295518 4224 295524 4236
rect 295576 4224 295582 4276
rect 88812 4168 89208 4196
rect 41874 4088 41880 4140
rect 41932 4128 41938 4140
rect 83458 4128 83464 4140
rect 41932 4100 83464 4128
rect 41932 4088 41938 4100
rect 83458 4088 83464 4100
rect 83516 4088 83522 4140
rect 85666 4088 85672 4140
rect 85724 4128 85730 4140
rect 88812 4128 88840 4168
rect 85724 4100 88840 4128
rect 88889 4131 88947 4137
rect 85724 4088 85730 4100
rect 88889 4097 88901 4131
rect 88935 4128 88947 4131
rect 89180 4128 89208 4168
rect 193214 4156 193220 4208
rect 193272 4196 193278 4208
rect 195238 4196 195244 4208
rect 193272 4168 195244 4196
rect 193272 4156 193278 4168
rect 195238 4156 195244 4168
rect 195296 4156 195302 4208
rect 225138 4156 225144 4208
rect 225196 4196 225202 4208
rect 228358 4196 228364 4208
rect 225196 4168 228364 4196
rect 225196 4156 225202 4168
rect 228358 4156 228364 4168
rect 228416 4156 228422 4208
rect 234522 4156 234528 4208
rect 234580 4196 234586 4208
rect 235810 4196 235816 4208
rect 234580 4168 235816 4196
rect 234580 4156 234586 4168
rect 235810 4156 235816 4168
rect 235868 4156 235874 4208
rect 280706 4156 280712 4208
rect 280764 4196 280770 4208
rect 285674 4196 285680 4208
rect 280764 4168 285680 4196
rect 280764 4156 280770 4168
rect 285674 4156 285680 4168
rect 285732 4156 285738 4208
rect 289078 4156 289084 4208
rect 289136 4196 289142 4208
rect 294874 4196 294880 4208
rect 289136 4168 294880 4196
rect 289136 4156 289142 4168
rect 294874 4156 294880 4168
rect 294932 4156 294938 4208
rect 497458 4156 497464 4208
rect 497516 4196 497522 4208
rect 498194 4196 498200 4208
rect 497516 4168 498200 4196
rect 497516 4156 497522 4168
rect 498194 4156 498200 4168
rect 498252 4156 498258 4208
rect 499574 4156 499580 4208
rect 499632 4196 499638 4208
rect 500586 4196 500592 4208
rect 499632 4168 500592 4196
rect 499632 4156 499638 4168
rect 500586 4156 500592 4168
rect 500644 4156 500650 4208
rect 522298 4156 522304 4208
rect 522356 4196 522362 4208
rect 523034 4196 523040 4208
rect 522356 4168 523040 4196
rect 522356 4156 522362 4168
rect 523034 4156 523040 4168
rect 523092 4156 523098 4208
rect 243170 4128 243176 4140
rect 88935 4100 89116 4128
rect 89180 4100 243176 4128
rect 88935 4097 88947 4100
rect 88889 4091 88947 4097
rect 60826 4020 60832 4072
rect 60884 4060 60890 4072
rect 65426 4060 65432 4072
rect 60884 4032 65432 4060
rect 60884 4020 60890 4032
rect 65426 4020 65432 4032
rect 65484 4020 65490 4072
rect 78582 4020 78588 4072
rect 78640 4060 78646 4072
rect 89088 4060 89116 4100
rect 243170 4088 243176 4100
rect 243228 4088 243234 4140
rect 257062 4088 257068 4140
rect 257120 4128 257126 4140
rect 260098 4128 260104 4140
rect 257120 4100 260104 4128
rect 257120 4088 257126 4100
rect 260098 4088 260104 4100
rect 260156 4088 260162 4140
rect 281350 4088 281356 4140
rect 281408 4128 281414 4140
rect 440326 4128 440332 4140
rect 281408 4100 440332 4128
rect 281408 4088 281414 4100
rect 440326 4088 440332 4100
rect 440384 4088 440390 4140
rect 453298 4088 453304 4140
rect 453356 4128 453362 4140
rect 560846 4128 560852 4140
rect 453356 4100 560852 4128
rect 453356 4088 453362 4100
rect 560846 4088 560852 4100
rect 560904 4088 560910 4140
rect 242986 4060 242992 4072
rect 78640 4032 89024 4060
rect 89088 4032 242992 4060
rect 78640 4020 78646 4032
rect 52546 3952 52552 4004
rect 52604 3992 52610 4004
rect 57238 3992 57244 4004
rect 52604 3964 57244 3992
rect 52604 3952 52610 3964
rect 57238 3952 57244 3964
rect 57296 3952 57302 4004
rect 82078 3952 82084 4004
rect 82136 3992 82142 4004
rect 88889 3995 88947 4001
rect 88889 3992 88901 3995
rect 82136 3964 88901 3992
rect 82136 3952 82142 3964
rect 88889 3961 88901 3964
rect 88935 3961 88947 3995
rect 88996 3992 89024 4032
rect 242986 4020 242992 4032
rect 243044 4020 243050 4072
rect 251174 4020 251180 4072
rect 251232 4060 251238 4072
rect 259914 4060 259920 4072
rect 251232 4032 259920 4060
rect 251232 4020 251238 4032
rect 259914 4020 259920 4032
rect 259972 4020 259978 4072
rect 281258 4020 281264 4072
rect 281316 4060 281322 4072
rect 436833 4063 436891 4069
rect 436833 4060 436845 4063
rect 281316 4032 436845 4060
rect 281316 4020 281322 4032
rect 436833 4029 436845 4032
rect 436879 4029 436891 4063
rect 436833 4023 436891 4029
rect 443638 4020 443644 4072
rect 443696 4060 443702 4072
rect 571518 4060 571524 4072
rect 443696 4032 571524 4060
rect 443696 4020 443702 4032
rect 571518 4020 571524 4032
rect 571576 4020 571582 4072
rect 243446 3992 243452 4004
rect 88996 3964 243452 3992
rect 88889 3955 88947 3961
rect 243446 3952 243452 3964
rect 243504 3952 243510 4004
rect 281166 3952 281172 4004
rect 281224 3992 281230 4004
rect 447410 3992 447416 4004
rect 281224 3964 447416 3992
rect 281224 3952 281230 3964
rect 447410 3952 447416 3964
rect 447468 3952 447474 4004
rect 450078 3992 450084 4004
rect 447704 3964 450084 3992
rect 44266 3884 44272 3936
rect 44324 3924 44330 3936
rect 50338 3924 50344 3936
rect 44324 3896 50344 3924
rect 44324 3884 44330 3896
rect 50338 3884 50344 3896
rect 50396 3884 50402 3936
rect 64322 3884 64328 3936
rect 64380 3924 64386 3936
rect 68370 3924 68376 3936
rect 64380 3896 68376 3924
rect 64380 3884 64386 3896
rect 68370 3884 68376 3896
rect 68428 3884 68434 3936
rect 74994 3884 75000 3936
rect 75052 3924 75058 3936
rect 241974 3924 241980 3936
rect 75052 3896 241980 3924
rect 75052 3884 75058 3896
rect 241974 3884 241980 3896
rect 242032 3884 242038 3936
rect 248782 3884 248788 3936
rect 248840 3924 248846 3936
rect 260190 3924 260196 3936
rect 248840 3896 260196 3924
rect 248840 3884 248846 3896
rect 260190 3884 260196 3896
rect 260248 3884 260254 3936
rect 281442 3884 281448 3936
rect 281500 3924 281506 3936
rect 447704 3924 447732 3964
rect 450078 3952 450084 3964
rect 450136 3952 450142 4004
rect 450538 3952 450544 4004
rect 450596 3992 450602 4004
rect 456061 3995 456119 4001
rect 450596 3964 452700 3992
rect 450596 3952 450602 3964
rect 281500 3896 447732 3924
rect 281500 3884 281506 3896
rect 447778 3884 447784 3936
rect 447836 3924 447842 3936
rect 452672 3924 452700 3964
rect 456061 3961 456073 3995
rect 456107 3992 456119 3995
rect 568022 3992 568028 4004
rect 456107 3964 568028 3992
rect 456107 3961 456119 3964
rect 456061 3955 456119 3961
rect 568022 3952 568028 3964
rect 568080 3952 568086 4004
rect 564434 3924 564440 3936
rect 447836 3896 452608 3924
rect 452672 3896 564440 3924
rect 447836 3884 447842 3896
rect 23014 3816 23020 3868
rect 23072 3856 23078 3868
rect 43438 3856 43444 3868
rect 23072 3828 43444 3856
rect 23072 3816 23078 3828
rect 43438 3816 43444 3828
rect 43496 3816 43502 3868
rect 46658 3816 46664 3868
rect 46716 3856 46722 3868
rect 239122 3856 239128 3868
rect 46716 3828 239128 3856
rect 46716 3816 46722 3828
rect 239122 3816 239128 3828
rect 239180 3816 239186 3868
rect 282822 3816 282828 3868
rect 282880 3856 282886 3868
rect 452580 3856 452608 3896
rect 564434 3884 564440 3896
rect 564492 3884 564498 3936
rect 456061 3859 456119 3865
rect 456061 3856 456073 3859
rect 282880 3828 452516 3856
rect 452580 3828 456073 3856
rect 282880 3816 282886 3828
rect 18230 3748 18236 3800
rect 18288 3788 18294 3800
rect 39390 3788 39396 3800
rect 18288 3760 39396 3788
rect 18288 3748 18294 3760
rect 39390 3748 39396 3760
rect 39448 3748 39454 3800
rect 43070 3748 43076 3800
rect 43128 3788 43134 3800
rect 233973 3791 234031 3797
rect 43128 3760 233924 3788
rect 43128 3748 43134 3760
rect 39574 3680 39580 3732
rect 39632 3720 39638 3732
rect 233896 3720 233924 3760
rect 233973 3757 233985 3791
rect 234019 3788 234031 3791
rect 238018 3788 238024 3800
rect 234019 3760 238024 3788
rect 234019 3757 234031 3760
rect 233973 3751 234031 3757
rect 238018 3748 238024 3760
rect 238076 3748 238082 3800
rect 255866 3748 255872 3800
rect 255924 3788 255930 3800
rect 260926 3788 260932 3800
rect 255924 3760 260932 3788
rect 255924 3748 255930 3760
rect 260926 3748 260932 3760
rect 260984 3748 260990 3800
rect 282638 3748 282644 3800
rect 282696 3788 282702 3800
rect 452381 3791 452439 3797
rect 452381 3788 452393 3791
rect 282696 3760 452393 3788
rect 282696 3748 282702 3760
rect 452381 3757 452393 3760
rect 452427 3757 452439 3791
rect 452488 3788 452516 3828
rect 456061 3825 456073 3828
rect 456107 3825 456119 3859
rect 550266 3856 550272 3868
rect 456061 3819 456119 3825
rect 456168 3828 550272 3856
rect 454494 3788 454500 3800
rect 452488 3760 454500 3788
rect 452381 3751 452439 3757
rect 454494 3748 454500 3760
rect 454552 3748 454558 3800
rect 454678 3748 454684 3800
rect 454736 3788 454742 3800
rect 456168 3788 456196 3828
rect 550266 3816 550272 3828
rect 550324 3816 550330 3868
rect 454736 3760 456196 3788
rect 454736 3748 454742 3760
rect 457438 3748 457444 3800
rect 457496 3788 457502 3800
rect 546678 3788 546684 3800
rect 457496 3760 546684 3788
rect 457496 3748 457502 3760
rect 546678 3748 546684 3760
rect 546736 3748 546742 3800
rect 239214 3720 239220 3732
rect 39632 3692 233832 3720
rect 233896 3692 239220 3720
rect 39632 3680 39638 3692
rect 32306 3612 32312 3664
rect 32364 3652 32370 3664
rect 32364 3624 35894 3652
rect 32364 3612 32370 3624
rect 27706 3544 27712 3596
rect 27764 3584 27770 3596
rect 28902 3584 28908 3596
rect 27764 3556 28908 3584
rect 27764 3544 27770 3556
rect 28902 3544 28908 3556
rect 28960 3544 28966 3596
rect 31294 3544 31300 3596
rect 31352 3584 31358 3596
rect 32490 3584 32496 3596
rect 31352 3556 32496 3584
rect 31352 3544 31358 3556
rect 32490 3544 32496 3556
rect 32548 3544 32554 3596
rect 33594 3544 33600 3596
rect 33652 3584 33658 3596
rect 34422 3584 34428 3596
rect 33652 3556 34428 3584
rect 33652 3544 33658 3556
rect 34422 3544 34428 3556
rect 34480 3544 34486 3596
rect 35866 3584 35894 3624
rect 35986 3612 35992 3664
rect 36044 3652 36050 3664
rect 233804 3652 233832 3692
rect 239214 3680 239220 3692
rect 239272 3680 239278 3732
rect 254670 3680 254676 3732
rect 254728 3720 254734 3732
rect 261202 3720 261208 3732
rect 254728 3692 261208 3720
rect 254728 3680 254734 3692
rect 261202 3680 261208 3692
rect 261260 3680 261266 3732
rect 282730 3680 282736 3732
rect 282788 3720 282794 3732
rect 461578 3720 461584 3732
rect 282788 3692 461584 3720
rect 282788 3680 282794 3692
rect 461578 3680 461584 3692
rect 461636 3680 461642 3732
rect 461670 3680 461676 3732
rect 461728 3720 461734 3732
rect 461728 3692 528554 3720
rect 461728 3680 461734 3692
rect 239398 3652 239404 3664
rect 36044 3624 233464 3652
rect 233804 3624 239404 3652
rect 36044 3612 36050 3624
rect 233329 3587 233387 3593
rect 233329 3584 233341 3587
rect 35866 3556 233341 3584
rect 233329 3553 233341 3556
rect 233375 3553 233387 3587
rect 233436 3584 233464 3624
rect 239398 3612 239404 3624
rect 239456 3612 239462 3664
rect 282546 3612 282552 3664
rect 282604 3652 282610 3664
rect 465166 3652 465172 3664
rect 282604 3624 465172 3652
rect 282604 3612 282610 3624
rect 465166 3612 465172 3624
rect 465224 3612 465230 3664
rect 468662 3652 468668 3664
rect 468404 3624 468668 3652
rect 237834 3584 237840 3596
rect 233436 3556 237840 3584
rect 233329 3547 233387 3553
rect 237834 3544 237840 3556
rect 237892 3544 237898 3596
rect 252370 3544 252376 3596
rect 252428 3584 252434 3596
rect 261018 3584 261024 3596
rect 252428 3556 261024 3584
rect 252428 3544 252434 3556
rect 261018 3544 261024 3556
rect 261076 3544 261082 3596
rect 263410 3544 263416 3596
rect 263468 3584 263474 3596
rect 266538 3584 266544 3596
rect 263468 3556 266544 3584
rect 263468 3544 263474 3556
rect 266538 3544 266544 3556
rect 266596 3544 266602 3596
rect 283742 3544 283748 3596
rect 283800 3584 283806 3596
rect 468404 3584 468432 3624
rect 468662 3612 468668 3624
rect 468720 3612 468726 3664
rect 528526 3652 528554 3692
rect 539594 3652 539600 3664
rect 528526 3624 539600 3652
rect 539594 3612 539600 3624
rect 539652 3612 539658 3664
rect 283800 3556 468432 3584
rect 283800 3544 283806 3556
rect 468478 3544 468484 3596
rect 468536 3584 468542 3596
rect 469858 3584 469864 3596
rect 468536 3556 469864 3584
rect 468536 3544 468542 3556
rect 469858 3544 469864 3556
rect 469916 3544 469922 3596
rect 514754 3544 514760 3596
rect 514812 3584 514818 3596
rect 515950 3584 515956 3596
rect 514812 3556 515956 3584
rect 514812 3544 514818 3556
rect 515950 3544 515956 3556
rect 516008 3544 516014 3596
rect 524414 3544 524420 3596
rect 524472 3584 524478 3596
rect 525426 3584 525432 3596
rect 524472 3556 525432 3584
rect 524472 3544 524478 3556
rect 525426 3544 525432 3556
rect 525484 3544 525490 3596
rect 17034 3476 17040 3528
rect 17092 3516 17098 3528
rect 17862 3516 17868 3528
rect 17092 3488 17868 3516
rect 17092 3476 17098 3488
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 25314 3476 25320 3528
rect 25372 3516 25378 3528
rect 25372 3488 229784 3516
rect 25372 3476 25378 3488
rect 13538 3408 13544 3460
rect 13596 3448 13602 3460
rect 22738 3448 22744 3460
rect 13596 3420 22744 3448
rect 13596 3408 13602 3420
rect 22738 3408 22744 3420
rect 22796 3408 22802 3460
rect 24210 3408 24216 3460
rect 24268 3448 24274 3460
rect 229281 3451 229339 3457
rect 229281 3448 229293 3451
rect 24268 3420 229293 3448
rect 24268 3408 24274 3420
rect 229281 3417 229293 3420
rect 229327 3417 229339 3451
rect 229756 3448 229784 3488
rect 229830 3476 229836 3528
rect 229888 3516 229894 3528
rect 230382 3516 230388 3528
rect 229888 3488 230388 3516
rect 229888 3476 229894 3488
rect 230382 3476 230388 3488
rect 230440 3476 230446 3528
rect 232222 3476 232228 3528
rect 232280 3516 232286 3528
rect 233142 3516 233148 3528
rect 232280 3488 233148 3516
rect 232280 3476 232286 3488
rect 233142 3476 233148 3488
rect 233200 3476 233206 3528
rect 233418 3476 233424 3528
rect 233476 3516 233482 3528
rect 234430 3516 234436 3528
rect 233476 3488 234436 3516
rect 233476 3476 233482 3488
rect 234430 3476 234436 3488
rect 234488 3476 234494 3528
rect 259454 3476 259460 3528
rect 259512 3516 259518 3528
rect 261110 3516 261116 3528
rect 259512 3488 261116 3516
rect 259512 3476 259518 3488
rect 261110 3476 261116 3488
rect 261168 3476 261174 3528
rect 262122 3476 262128 3528
rect 262180 3516 262186 3528
rect 262950 3516 262956 3528
rect 262180 3488 262956 3516
rect 262180 3476 262186 3488
rect 262950 3476 262956 3488
rect 263008 3476 263014 3528
rect 264238 3476 264244 3528
rect 264296 3516 264302 3528
rect 265342 3516 265348 3528
rect 264296 3488 265348 3516
rect 264296 3476 264302 3488
rect 265342 3476 265348 3488
rect 265400 3476 265406 3528
rect 283926 3476 283932 3528
rect 283984 3516 283990 3528
rect 472250 3516 472256 3528
rect 283984 3488 472256 3516
rect 283984 3476 283990 3488
rect 472250 3476 472256 3488
rect 472308 3476 472314 3528
rect 475746 3516 475752 3528
rect 472544 3488 475752 3516
rect 237650 3448 237656 3460
rect 229756 3420 237656 3448
rect 229281 3411 229339 3417
rect 237650 3408 237656 3420
rect 237708 3408 237714 3460
rect 245194 3408 245200 3460
rect 245252 3448 245258 3460
rect 257338 3448 257344 3460
rect 245252 3420 257344 3448
rect 245252 3408 245258 3420
rect 257338 3408 257344 3420
rect 257396 3408 257402 3460
rect 262858 3408 262864 3460
rect 262916 3448 262922 3460
rect 264146 3448 264152 3460
rect 262916 3420 264152 3448
rect 262916 3408 262922 3420
rect 264146 3408 264152 3420
rect 264204 3408 264210 3460
rect 284018 3408 284024 3460
rect 284076 3448 284082 3460
rect 472544 3448 472572 3488
rect 475746 3476 475752 3488
rect 475804 3476 475810 3528
rect 510062 3476 510068 3528
rect 510120 3516 510126 3528
rect 510706 3516 510712 3528
rect 510120 3488 510712 3516
rect 510120 3476 510126 3488
rect 510706 3476 510712 3488
rect 510764 3476 510770 3528
rect 512638 3476 512644 3528
rect 512696 3516 512702 3528
rect 513558 3516 513564 3528
rect 512696 3488 513564 3516
rect 512696 3476 512702 3488
rect 513558 3476 513564 3488
rect 513616 3476 513622 3528
rect 519538 3476 519544 3528
rect 519596 3516 519602 3528
rect 521838 3516 521844 3528
rect 519596 3488 521844 3516
rect 519596 3476 519602 3488
rect 521838 3476 521844 3488
rect 521896 3476 521902 3528
rect 530578 3476 530584 3528
rect 530636 3516 530642 3528
rect 531314 3516 531320 3528
rect 530636 3488 531320 3516
rect 530636 3476 530642 3488
rect 531314 3476 531320 3488
rect 531372 3476 531378 3528
rect 534902 3476 534908 3528
rect 534960 3516 534966 3528
rect 535454 3516 535460 3528
rect 534960 3488 535460 3516
rect 534960 3476 534966 3488
rect 535454 3476 535460 3488
rect 535512 3476 535518 3528
rect 541986 3476 541992 3528
rect 542044 3516 542050 3528
rect 542446 3516 542452 3528
rect 542044 3488 542452 3516
rect 542044 3476 542050 3488
rect 542446 3476 542452 3488
rect 542504 3476 542510 3528
rect 545482 3476 545488 3528
rect 545540 3516 545546 3528
rect 546494 3516 546500 3528
rect 545540 3488 546500 3516
rect 545540 3476 545546 3488
rect 546494 3476 546500 3488
rect 546552 3476 546558 3528
rect 551278 3476 551284 3528
rect 551336 3516 551342 3528
rect 552658 3516 552664 3528
rect 551336 3488 552664 3516
rect 551336 3476 551342 3488
rect 552658 3476 552664 3488
rect 552716 3476 552722 3528
rect 559742 3476 559748 3528
rect 559800 3516 559806 3528
rect 560294 3516 560300 3528
rect 559800 3488 560300 3516
rect 559800 3476 559806 3488
rect 560294 3476 560300 3488
rect 560352 3476 560358 3528
rect 284076 3420 472572 3448
rect 284076 3408 284082 3420
rect 472618 3408 472624 3460
rect 472676 3448 472682 3460
rect 473446 3448 473452 3460
rect 472676 3420 473452 3448
rect 472676 3408 472682 3420
rect 473446 3408 473452 3420
rect 473504 3408 473510 3460
rect 483750 3408 483756 3460
rect 483808 3448 483814 3460
rect 553762 3448 553768 3460
rect 483808 3420 553768 3448
rect 483808 3408 483814 3420
rect 553762 3408 553768 3420
rect 553820 3408 553826 3460
rect 566550 3408 566556 3460
rect 566608 3448 566614 3460
rect 572714 3448 572720 3460
rect 566608 3420 572720 3448
rect 566608 3408 566614 3420
rect 572714 3408 572720 3420
rect 572772 3408 572778 3460
rect 26510 3340 26516 3392
rect 26568 3380 26574 3392
rect 29638 3380 29644 3392
rect 26568 3352 29644 3380
rect 26568 3340 26574 3352
rect 29638 3340 29644 3352
rect 29696 3340 29702 3392
rect 30098 3340 30104 3392
rect 30156 3380 30162 3392
rect 32398 3380 32404 3392
rect 30156 3352 32404 3380
rect 30156 3340 30162 3352
rect 32398 3340 32404 3352
rect 32456 3340 32462 3392
rect 34790 3340 34796 3392
rect 34848 3380 34854 3392
rect 35802 3380 35808 3392
rect 34848 3352 35808 3380
rect 34848 3340 34854 3352
rect 35802 3340 35808 3352
rect 35860 3340 35866 3392
rect 38378 3340 38384 3392
rect 38436 3380 38442 3392
rect 39298 3380 39304 3392
rect 38436 3352 39304 3380
rect 38436 3340 38442 3352
rect 39298 3340 39304 3352
rect 39356 3340 39362 3392
rect 40678 3340 40684 3392
rect 40736 3380 40742 3392
rect 41322 3380 41328 3392
rect 40736 3352 41328 3380
rect 40736 3340 40742 3352
rect 41322 3340 41328 3352
rect 41380 3340 41386 3392
rect 50154 3340 50160 3392
rect 50212 3380 50218 3392
rect 50982 3380 50988 3392
rect 50212 3352 50988 3380
rect 50212 3340 50218 3352
rect 50982 3340 50988 3352
rect 51040 3340 51046 3392
rect 51350 3340 51356 3392
rect 51408 3380 51414 3392
rect 52362 3380 52368 3392
rect 51408 3352 52368 3380
rect 51408 3340 51414 3352
rect 52362 3340 52368 3352
rect 52420 3340 52426 3392
rect 56042 3340 56048 3392
rect 56100 3380 56106 3392
rect 57330 3380 57336 3392
rect 56100 3352 57336 3380
rect 56100 3340 56106 3352
rect 57330 3340 57336 3352
rect 57388 3340 57394 3392
rect 58434 3340 58440 3392
rect 58492 3380 58498 3392
rect 59262 3380 59268 3392
rect 58492 3352 59268 3380
rect 58492 3340 58498 3352
rect 59262 3340 59268 3352
rect 59320 3340 59326 3392
rect 59630 3340 59636 3392
rect 59688 3380 59694 3392
rect 61378 3380 61384 3392
rect 59688 3352 61384 3380
rect 59688 3340 59694 3352
rect 61378 3340 61384 3352
rect 61436 3340 61442 3392
rect 65518 3340 65524 3392
rect 65576 3380 65582 3392
rect 66162 3380 66168 3392
rect 65576 3352 66168 3380
rect 65576 3340 65582 3352
rect 66162 3340 66168 3352
rect 66220 3340 66226 3392
rect 66714 3340 66720 3392
rect 66772 3380 66778 3392
rect 68278 3380 68284 3392
rect 66772 3352 68284 3380
rect 66772 3340 66778 3352
rect 68278 3340 68284 3352
rect 68336 3340 68342 3392
rect 69106 3340 69112 3392
rect 69164 3380 69170 3392
rect 70210 3380 70216 3392
rect 69164 3352 70216 3380
rect 69164 3340 69170 3352
rect 70210 3340 70216 3352
rect 70268 3340 70274 3392
rect 70302 3340 70308 3392
rect 70360 3380 70366 3392
rect 71038 3380 71044 3392
rect 70360 3352 71044 3380
rect 70360 3340 70366 3352
rect 71038 3340 71044 3352
rect 71096 3340 71102 3392
rect 72602 3340 72608 3392
rect 72660 3380 72666 3392
rect 73062 3380 73068 3392
rect 72660 3352 73068 3380
rect 72660 3340 72666 3352
rect 73062 3340 73068 3352
rect 73120 3340 73126 3392
rect 76190 3340 76196 3392
rect 76248 3380 76254 3392
rect 77202 3380 77208 3392
rect 76248 3352 77208 3380
rect 76248 3340 76254 3352
rect 77202 3340 77208 3352
rect 77260 3340 77266 3392
rect 77386 3340 77392 3392
rect 77444 3380 77450 3392
rect 79318 3380 79324 3392
rect 77444 3352 79324 3380
rect 77444 3340 77450 3352
rect 79318 3340 79324 3352
rect 79376 3340 79382 3392
rect 80882 3340 80888 3392
rect 80940 3380 80946 3392
rect 81342 3380 81348 3392
rect 80940 3352 81348 3380
rect 80940 3340 80946 3352
rect 81342 3340 81348 3352
rect 81400 3340 81406 3392
rect 90358 3340 90364 3392
rect 90416 3380 90422 3392
rect 91002 3380 91008 3392
rect 90416 3352 91008 3380
rect 90416 3340 90422 3352
rect 91002 3340 91008 3352
rect 91060 3340 91066 3392
rect 91554 3340 91560 3392
rect 91612 3380 91618 3392
rect 93118 3380 93124 3392
rect 91612 3352 93124 3380
rect 91612 3340 91618 3352
rect 93118 3340 93124 3352
rect 93176 3340 93182 3392
rect 93946 3340 93952 3392
rect 94004 3380 94010 3392
rect 95050 3380 95056 3392
rect 94004 3352 95056 3380
rect 94004 3340 94010 3352
rect 95050 3340 95056 3352
rect 95108 3340 95114 3392
rect 97442 3340 97448 3392
rect 97500 3380 97506 3392
rect 97902 3380 97908 3392
rect 97500 3352 97908 3380
rect 97500 3340 97506 3352
rect 97902 3340 97908 3352
rect 97960 3340 97966 3392
rect 98638 3340 98644 3392
rect 98696 3380 98702 3392
rect 99282 3380 99288 3392
rect 98696 3352 99288 3380
rect 98696 3340 98702 3352
rect 99282 3340 99288 3352
rect 99340 3340 99346 3392
rect 101030 3340 101036 3392
rect 101088 3380 101094 3392
rect 102042 3380 102048 3392
rect 101088 3352 102048 3380
rect 101088 3340 101094 3352
rect 102042 3340 102048 3352
rect 102100 3340 102106 3392
rect 243078 3380 243084 3392
rect 102152 3352 243084 3380
rect 67910 3272 67916 3324
rect 67968 3312 67974 3324
rect 69658 3312 69664 3324
rect 67968 3284 69664 3312
rect 67968 3272 67974 3284
rect 69658 3272 69664 3284
rect 69716 3272 69722 3324
rect 87966 3272 87972 3324
rect 88024 3312 88030 3324
rect 88978 3312 88984 3324
rect 88024 3284 88984 3312
rect 88024 3272 88030 3284
rect 88978 3272 88984 3284
rect 89036 3272 89042 3324
rect 11146 3204 11152 3256
rect 11204 3244 11210 3256
rect 14458 3244 14464 3256
rect 11204 3216 14464 3244
rect 11204 3204 11210 3216
rect 14458 3204 14464 3216
rect 14516 3204 14522 3256
rect 57238 3204 57244 3256
rect 57296 3244 57302 3256
rect 58618 3244 58624 3256
rect 57296 3216 58624 3244
rect 57296 3204 57302 3216
rect 58618 3204 58624 3216
rect 58676 3204 58682 3256
rect 89162 3204 89168 3256
rect 89220 3244 89226 3256
rect 102152 3244 102180 3352
rect 243078 3340 243084 3352
rect 243136 3340 243142 3392
rect 279970 3340 279976 3392
rect 280028 3380 280034 3392
rect 280028 3352 431954 3380
rect 280028 3340 280034 3352
rect 102229 3315 102287 3321
rect 102229 3281 102241 3315
rect 102275 3312 102287 3315
rect 244550 3312 244556 3324
rect 102275 3284 244556 3312
rect 102275 3281 102287 3284
rect 102229 3275 102287 3281
rect 244550 3272 244556 3284
rect 244608 3272 244614 3324
rect 279786 3272 279792 3324
rect 279844 3312 279850 3324
rect 279844 3284 425652 3312
rect 279844 3272 279850 3284
rect 244734 3244 244740 3256
rect 89220 3216 102180 3244
rect 102244 3216 244740 3244
rect 89220 3204 89226 3216
rect 48958 3068 48964 3120
rect 49016 3108 49022 3120
rect 53098 3108 53104 3120
rect 49016 3080 53104 3108
rect 49016 3068 49022 3080
rect 53098 3068 53104 3080
rect 53156 3068 53162 3120
rect 96246 3068 96252 3120
rect 96304 3108 96310 3120
rect 102244 3108 102272 3216
rect 244734 3204 244740 3216
rect 244792 3204 244798 3256
rect 279878 3204 279884 3256
rect 279936 3244 279942 3256
rect 425624 3244 425652 3284
rect 425698 3272 425704 3324
rect 425756 3312 425762 3324
rect 427262 3312 427268 3324
rect 425756 3284 427268 3312
rect 425756 3272 425762 3284
rect 427262 3272 427268 3284
rect 427320 3272 427326 3324
rect 431926 3312 431954 3352
rect 432598 3340 432604 3392
rect 432656 3380 432662 3392
rect 434438 3380 434444 3392
rect 432656 3352 434444 3380
rect 432656 3340 432662 3352
rect 434438 3340 434444 3352
rect 434496 3340 434502 3392
rect 436738 3340 436744 3392
rect 436796 3380 436802 3392
rect 437934 3380 437940 3392
rect 436796 3352 437940 3380
rect 436796 3340 436802 3352
rect 437934 3340 437940 3352
rect 437992 3340 437998 3392
rect 448514 3340 448520 3392
rect 448572 3380 448578 3392
rect 449802 3380 449808 3392
rect 448572 3352 449808 3380
rect 448572 3340 448578 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 452381 3383 452439 3389
rect 452381 3349 452393 3383
rect 452427 3380 452439 3383
rect 458082 3380 458088 3392
rect 452427 3352 458088 3380
rect 452427 3349 452439 3352
rect 452381 3343 452439 3349
rect 458082 3340 458088 3352
rect 458140 3340 458146 3392
rect 464338 3340 464344 3392
rect 464396 3380 464402 3392
rect 536098 3380 536104 3392
rect 464396 3352 536104 3380
rect 464396 3340 464402 3352
rect 536098 3340 536104 3352
rect 536156 3340 536162 3392
rect 436833 3315 436891 3321
rect 431926 3284 436784 3312
rect 436756 3256 436784 3284
rect 436833 3281 436845 3315
rect 436879 3312 436891 3315
rect 443822 3312 443828 3324
rect 436879 3284 443828 3312
rect 436879 3281 436891 3284
rect 436833 3275 436891 3281
rect 443822 3272 443828 3284
rect 443880 3272 443886 3324
rect 433242 3244 433248 3256
rect 279936 3216 425468 3244
rect 425624 3216 433248 3244
rect 279936 3204 279942 3216
rect 102321 3179 102379 3185
rect 102321 3145 102333 3179
rect 102367 3176 102379 3179
rect 244826 3176 244832 3188
rect 102367 3148 244832 3176
rect 102367 3145 102379 3148
rect 102321 3139 102379 3145
rect 244826 3136 244832 3148
rect 244884 3136 244890 3188
rect 258258 3136 258264 3188
rect 258316 3176 258322 3188
rect 261294 3176 261300 3188
rect 258316 3148 261300 3176
rect 258316 3136 258322 3148
rect 261294 3136 261300 3148
rect 261352 3136 261358 3188
rect 263502 3136 263508 3188
rect 263560 3176 263566 3188
rect 270034 3176 270040 3188
rect 263560 3148 270040 3176
rect 263560 3136 263566 3148
rect 270034 3136 270040 3148
rect 270092 3136 270098 3188
rect 279602 3136 279608 3188
rect 279660 3176 279666 3188
rect 279660 3148 413324 3176
rect 279660 3136 279666 3148
rect 96304 3080 102272 3108
rect 96304 3068 96310 3080
rect 103330 3068 103336 3120
rect 103388 3108 103394 3120
rect 245102 3108 245108 3120
rect 103388 3080 245108 3108
rect 103388 3068 103394 3080
rect 245102 3068 245108 3080
rect 245160 3068 245166 3120
rect 278130 3068 278136 3120
rect 278188 3108 278194 3120
rect 413296 3108 413324 3148
rect 414658 3136 414664 3188
rect 414716 3176 414722 3188
rect 416682 3176 416688 3188
rect 414716 3148 416688 3176
rect 414716 3136 414722 3148
rect 416682 3136 416688 3148
rect 416740 3136 416746 3188
rect 278188 3080 409460 3108
rect 413296 3080 418154 3108
rect 278188 3068 278194 3080
rect 19426 3000 19432 3052
rect 19484 3040 19490 3052
rect 25498 3040 25504 3052
rect 19484 3012 25504 3040
rect 19484 3000 19490 3012
rect 25498 3000 25504 3012
rect 25556 3000 25562 3052
rect 92750 3000 92756 3052
rect 92808 3040 92814 3052
rect 102229 3043 102287 3049
rect 102229 3040 102241 3043
rect 92808 3012 102241 3040
rect 92808 3000 92814 3012
rect 102229 3009 102241 3012
rect 102275 3009 102287 3043
rect 102229 3003 102287 3009
rect 105722 3000 105728 3052
rect 105780 3040 105786 3052
rect 106182 3040 106188 3052
rect 105780 3012 106188 3040
rect 105780 3000 105786 3012
rect 106182 3000 106188 3012
rect 106240 3000 106246 3052
rect 106918 3000 106924 3052
rect 106976 3040 106982 3052
rect 107562 3040 107568 3052
rect 106976 3012 107568 3040
rect 106976 3000 106982 3012
rect 107562 3000 107568 3012
rect 107620 3000 107626 3052
rect 108114 3000 108120 3052
rect 108172 3040 108178 3052
rect 108942 3040 108948 3052
rect 108172 3012 108948 3040
rect 108172 3000 108178 3012
rect 108942 3000 108948 3012
rect 109000 3000 109006 3052
rect 109310 3000 109316 3052
rect 109368 3040 109374 3052
rect 111058 3040 111064 3052
rect 109368 3012 111064 3040
rect 109368 3000 109374 3012
rect 111058 3000 111064 3012
rect 111116 3000 111122 3052
rect 111150 3000 111156 3052
rect 111208 3040 111214 3052
rect 246206 3040 246212 3052
rect 111208 3012 246212 3040
rect 111208 3000 111214 3012
rect 246206 3000 246212 3012
rect 246264 3000 246270 3052
rect 263318 3000 263324 3052
rect 263376 3040 263382 3052
rect 268838 3040 268844 3052
rect 263376 3012 268844 3040
rect 263376 3000 263382 3012
rect 268838 3000 268844 3012
rect 268896 3000 268902 3052
rect 277946 3000 277952 3052
rect 278004 3040 278010 3052
rect 278004 3012 409368 3040
rect 278004 3000 278010 3012
rect 73798 2932 73804 2984
rect 73856 2972 73862 2984
rect 75178 2972 75184 2984
rect 73856 2944 75184 2972
rect 73856 2932 73862 2944
rect 75178 2932 75184 2944
rect 75236 2932 75242 2984
rect 115106 2972 115112 2984
rect 84166 2944 115112 2972
rect 71498 2864 71504 2916
rect 71556 2904 71562 2916
rect 84166 2904 84194 2944
rect 115106 2932 115112 2944
rect 115164 2932 115170 2984
rect 115198 2932 115204 2984
rect 115256 2972 115262 2984
rect 115842 2972 115848 2984
rect 115256 2944 115848 2972
rect 115256 2932 115262 2944
rect 115842 2932 115848 2944
rect 115900 2932 115906 2984
rect 116394 2932 116400 2984
rect 116452 2972 116458 2984
rect 117222 2972 117228 2984
rect 116452 2944 117228 2972
rect 116452 2932 116458 2944
rect 117222 2932 117228 2944
rect 117280 2932 117286 2984
rect 118786 2932 118792 2984
rect 118844 2972 118850 2984
rect 119798 2972 119804 2984
rect 118844 2944 119804 2972
rect 118844 2932 118850 2944
rect 119798 2932 119804 2944
rect 119856 2932 119862 2984
rect 122098 2972 122104 2984
rect 119908 2944 122104 2972
rect 71556 2876 84194 2904
rect 71556 2864 71562 2876
rect 84470 2864 84476 2916
rect 84528 2904 84534 2916
rect 87598 2904 87604 2916
rect 84528 2876 87604 2904
rect 84528 2864 84534 2876
rect 87598 2864 87604 2876
rect 87656 2864 87662 2916
rect 99834 2864 99840 2916
rect 99892 2904 99898 2916
rect 102321 2907 102379 2913
rect 102321 2904 102333 2907
rect 99892 2876 102333 2904
rect 99892 2864 99898 2876
rect 102321 2873 102333 2876
rect 102367 2873 102379 2907
rect 102321 2867 102379 2873
rect 114002 2864 114008 2916
rect 114060 2904 114066 2916
rect 119908 2904 119936 2944
rect 122098 2932 122104 2944
rect 122156 2932 122162 2984
rect 122282 2932 122288 2984
rect 122340 2972 122346 2984
rect 122742 2972 122748 2984
rect 122340 2944 122748 2972
rect 122340 2932 122346 2944
rect 122742 2932 122748 2944
rect 122800 2932 122806 2984
rect 123478 2932 123484 2984
rect 123536 2972 123542 2984
rect 124122 2972 124128 2984
rect 123536 2944 124128 2972
rect 123536 2932 123542 2944
rect 124122 2932 124128 2944
rect 124180 2932 124186 2984
rect 124674 2932 124680 2984
rect 124732 2972 124738 2984
rect 125410 2972 125416 2984
rect 124732 2944 125416 2972
rect 124732 2932 124738 2944
rect 125410 2932 125416 2944
rect 125468 2932 125474 2984
rect 125870 2932 125876 2984
rect 125928 2972 125934 2984
rect 126882 2972 126888 2984
rect 125928 2944 126888 2972
rect 125928 2932 125934 2944
rect 126882 2932 126888 2944
rect 126940 2932 126946 2984
rect 126974 2932 126980 2984
rect 127032 2972 127038 2984
rect 128998 2972 129004 2984
rect 127032 2944 129004 2972
rect 127032 2932 127038 2944
rect 128998 2932 129004 2944
rect 129056 2932 129062 2984
rect 129093 2975 129151 2981
rect 129093 2941 129105 2975
rect 129139 2972 129151 2975
rect 246114 2972 246120 2984
rect 129139 2944 246120 2972
rect 129139 2941 129151 2944
rect 129093 2935 129151 2941
rect 246114 2932 246120 2944
rect 246172 2932 246178 2984
rect 278498 2932 278504 2984
rect 278556 2972 278562 2984
rect 409233 2975 409291 2981
rect 409233 2972 409245 2975
rect 278556 2944 409245 2972
rect 278556 2932 278562 2944
rect 409233 2941 409245 2944
rect 409279 2941 409291 2975
rect 409233 2935 409291 2941
rect 114060 2876 119936 2904
rect 114060 2864 114066 2876
rect 121086 2864 121092 2916
rect 121144 2904 121150 2916
rect 247494 2904 247500 2916
rect 121144 2876 129044 2904
rect 121144 2864 121150 2876
rect 110506 2796 110512 2848
rect 110564 2836 110570 2848
rect 111150 2836 111156 2848
rect 110564 2808 111156 2836
rect 110564 2796 110570 2808
rect 111150 2796 111156 2808
rect 111208 2796 111214 2848
rect 117590 2796 117596 2848
rect 117648 2836 117654 2848
rect 128909 2839 128967 2845
rect 128909 2836 128921 2839
rect 117648 2808 128921 2836
rect 117648 2796 117654 2808
rect 128909 2805 128921 2808
rect 128955 2805 128967 2839
rect 128909 2799 128967 2805
rect 129016 2768 129044 2876
rect 132466 2876 247500 2904
rect 132466 2836 132494 2876
rect 247494 2864 247500 2876
rect 247552 2864 247558 2916
rect 276750 2864 276756 2916
rect 276808 2904 276814 2916
rect 276808 2876 396672 2904
rect 276808 2864 276814 2876
rect 129200 2808 132494 2836
rect 129200 2768 129228 2808
rect 132954 2796 132960 2848
rect 133012 2836 133018 2848
rect 133782 2836 133788 2848
rect 133012 2808 133788 2836
rect 133012 2796 133018 2808
rect 133782 2796 133788 2808
rect 133840 2796 133846 2848
rect 134150 2796 134156 2848
rect 134208 2836 134214 2848
rect 135162 2836 135168 2848
rect 134208 2808 135168 2836
rect 134208 2796 134214 2808
rect 135162 2796 135168 2808
rect 135220 2796 135226 2848
rect 136450 2796 136456 2848
rect 136508 2836 136514 2848
rect 137278 2836 137284 2848
rect 136508 2808 137284 2836
rect 136508 2796 136514 2808
rect 137278 2796 137284 2808
rect 137336 2796 137342 2848
rect 140038 2796 140044 2848
rect 140096 2836 140102 2848
rect 140682 2836 140688 2848
rect 140096 2808 140688 2836
rect 140096 2796 140102 2808
rect 140682 2796 140688 2808
rect 140740 2796 140746 2848
rect 141234 2796 141240 2848
rect 141292 2836 141298 2848
rect 142062 2836 142068 2848
rect 141292 2808 142068 2836
rect 141292 2796 141298 2808
rect 142062 2796 142068 2808
rect 142120 2796 142126 2848
rect 143534 2796 143540 2848
rect 143592 2836 143598 2848
rect 144822 2836 144828 2848
rect 143592 2808 144828 2836
rect 143592 2796 143598 2808
rect 144822 2796 144828 2808
rect 144880 2796 144886 2848
rect 147122 2796 147128 2848
rect 147180 2836 147186 2848
rect 147582 2836 147588 2848
rect 147180 2808 147588 2836
rect 147180 2796 147186 2808
rect 147582 2796 147588 2808
rect 147640 2796 147646 2848
rect 148318 2796 148324 2848
rect 148376 2836 148382 2848
rect 148962 2836 148968 2848
rect 148376 2808 148968 2836
rect 148376 2796 148382 2808
rect 148962 2796 148968 2808
rect 149020 2796 149026 2848
rect 149514 2796 149520 2848
rect 149572 2836 149578 2848
rect 150342 2836 150348 2848
rect 149572 2808 150348 2836
rect 149572 2796 149578 2808
rect 150342 2796 150348 2808
rect 150400 2796 150406 2848
rect 150618 2796 150624 2848
rect 150676 2836 150682 2848
rect 151722 2836 151728 2848
rect 150676 2808 151728 2836
rect 150676 2796 150682 2808
rect 151722 2796 151728 2808
rect 151780 2796 151786 2848
rect 151814 2796 151820 2848
rect 151872 2836 151878 2848
rect 153102 2836 153108 2848
rect 151872 2808 153108 2836
rect 151872 2796 151878 2808
rect 153102 2796 153108 2808
rect 153160 2796 153166 2848
rect 154206 2796 154212 2848
rect 154264 2836 154270 2848
rect 155218 2836 155224 2848
rect 154264 2808 155224 2836
rect 154264 2796 154270 2808
rect 155218 2796 155224 2808
rect 155276 2796 155282 2848
rect 155402 2796 155408 2848
rect 155460 2836 155466 2848
rect 155862 2836 155868 2848
rect 155460 2808 155868 2836
rect 155460 2796 155466 2808
rect 155862 2796 155868 2808
rect 155920 2796 155926 2848
rect 156598 2796 156604 2848
rect 156656 2836 156662 2848
rect 157242 2836 157248 2848
rect 156656 2808 157248 2836
rect 156656 2796 156662 2808
rect 157242 2796 157248 2808
rect 157300 2796 157306 2848
rect 157794 2796 157800 2848
rect 157852 2836 157858 2848
rect 158622 2836 158628 2848
rect 157852 2808 158628 2836
rect 157852 2796 157858 2808
rect 158622 2796 158628 2808
rect 158680 2796 158686 2848
rect 164878 2796 164884 2848
rect 164936 2836 164942 2848
rect 165522 2836 165528 2848
rect 164936 2808 165528 2836
rect 164936 2796 164942 2808
rect 165522 2796 165528 2808
rect 165580 2796 165586 2848
rect 166074 2796 166080 2848
rect 166132 2836 166138 2848
rect 166902 2836 166908 2848
rect 166132 2808 166908 2836
rect 166132 2796 166138 2808
rect 166902 2796 166908 2808
rect 166960 2796 166966 2848
rect 168374 2796 168380 2848
rect 168432 2836 168438 2848
rect 169662 2836 169668 2848
rect 168432 2808 169668 2836
rect 168432 2796 168438 2808
rect 169662 2796 169668 2808
rect 169720 2796 169726 2848
rect 188522 2796 188528 2848
rect 188580 2836 188586 2848
rect 188982 2836 188988 2848
rect 188580 2808 188988 2836
rect 188580 2796 188586 2808
rect 188982 2796 188988 2808
rect 189040 2796 189046 2848
rect 190822 2796 190828 2848
rect 190880 2836 190886 2848
rect 191742 2836 191748 2848
rect 190880 2808 191748 2836
rect 190880 2796 190886 2808
rect 191742 2796 191748 2808
rect 191800 2796 191806 2848
rect 192018 2796 192024 2848
rect 192076 2836 192082 2848
rect 193122 2836 193128 2848
rect 192076 2808 193128 2836
rect 192076 2796 192082 2808
rect 193122 2796 193128 2808
rect 193180 2796 193186 2848
rect 197906 2796 197912 2848
rect 197964 2836 197970 2848
rect 198642 2836 198648 2848
rect 197964 2808 198648 2836
rect 197964 2796 197970 2808
rect 198642 2796 198648 2808
rect 198700 2796 198706 2848
rect 206186 2796 206192 2848
rect 206244 2836 206250 2848
rect 206922 2836 206928 2848
rect 206244 2808 206928 2836
rect 206244 2796 206250 2808
rect 206922 2796 206928 2808
rect 206980 2796 206986 2848
rect 209774 2796 209780 2848
rect 209832 2836 209838 2848
rect 210970 2836 210976 2848
rect 209832 2808 210976 2836
rect 209832 2796 209838 2808
rect 210970 2796 210976 2808
rect 211028 2796 211034 2848
rect 213362 2796 213368 2848
rect 213420 2836 213426 2848
rect 213822 2836 213828 2848
rect 213420 2808 213828 2836
rect 213420 2796 213426 2808
rect 213822 2796 213828 2808
rect 213880 2796 213886 2848
rect 214466 2796 214472 2848
rect 214524 2836 214530 2848
rect 215202 2836 215208 2848
rect 214524 2808 215208 2836
rect 214524 2796 214530 2808
rect 215202 2796 215208 2808
rect 215260 2796 215266 2848
rect 215662 2796 215668 2848
rect 215720 2836 215726 2848
rect 216582 2836 216588 2848
rect 215720 2808 216588 2836
rect 215720 2796 215726 2808
rect 216582 2796 216588 2808
rect 216640 2796 216646 2848
rect 216858 2796 216864 2848
rect 216916 2836 216922 2848
rect 217962 2836 217968 2848
rect 216916 2808 217968 2836
rect 216916 2796 216922 2808
rect 217962 2796 217968 2808
rect 218020 2796 218026 2848
rect 219250 2796 219256 2848
rect 219308 2836 219314 2848
rect 220078 2836 220084 2848
rect 219308 2808 220084 2836
rect 219308 2796 219314 2808
rect 220078 2796 220084 2808
rect 220136 2796 220142 2848
rect 222746 2796 222752 2848
rect 222804 2836 222810 2848
rect 223482 2836 223488 2848
rect 222804 2808 223488 2836
rect 222804 2796 222810 2808
rect 223482 2796 223488 2808
rect 223540 2796 223546 2848
rect 223942 2796 223948 2848
rect 224000 2836 224006 2848
rect 224862 2836 224868 2848
rect 224000 2808 224868 2836
rect 224000 2796 224006 2808
rect 224862 2796 224868 2808
rect 224920 2796 224926 2848
rect 226334 2796 226340 2848
rect 226392 2836 226398 2848
rect 227438 2836 227444 2848
rect 226392 2808 227444 2836
rect 226392 2796 226398 2808
rect 227438 2796 227444 2808
rect 227496 2796 227502 2848
rect 229281 2839 229339 2845
rect 229281 2805 229293 2839
rect 229327 2836 229339 2839
rect 237926 2836 237932 2848
rect 229327 2808 237932 2836
rect 229327 2805 229339 2808
rect 229281 2799 229339 2805
rect 237926 2796 237932 2808
rect 237984 2796 237990 2848
rect 300118 2796 300124 2848
rect 300176 2836 300182 2848
rect 301958 2836 301964 2848
rect 300176 2808 301964 2836
rect 300176 2796 300182 2808
rect 301958 2796 301964 2808
rect 302016 2796 302022 2848
rect 307018 2796 307024 2848
rect 307076 2836 307082 2848
rect 307938 2836 307944 2848
rect 307076 2808 307944 2836
rect 307076 2796 307082 2808
rect 307938 2796 307944 2808
rect 307996 2796 308002 2848
rect 313918 2796 313924 2848
rect 313976 2836 313982 2848
rect 315022 2836 315028 2848
rect 313976 2808 315028 2836
rect 313976 2796 313982 2808
rect 315022 2796 315028 2808
rect 315080 2796 315086 2848
rect 316034 2796 316040 2848
rect 316092 2836 316098 2848
rect 317322 2836 317328 2848
rect 316092 2808 317328 2836
rect 316092 2796 316098 2808
rect 317322 2796 317328 2808
rect 317380 2796 317386 2848
rect 331950 2796 331956 2848
rect 332008 2836 332014 2848
rect 332008 2808 332640 2836
rect 332008 2796 332014 2808
rect 129016 2740 129228 2768
rect 332612 2768 332640 2808
rect 332686 2796 332692 2848
rect 332744 2836 332750 2848
rect 333974 2836 333980 2848
rect 332744 2808 333980 2836
rect 332744 2796 332750 2808
rect 333974 2796 333980 2808
rect 334032 2796 334038 2848
rect 337470 2796 337476 2848
rect 337528 2836 337534 2848
rect 338114 2836 338120 2848
rect 337528 2808 338120 2836
rect 337528 2796 337534 2808
rect 338114 2796 338120 2808
rect 338172 2796 338178 2848
rect 342990 2796 342996 2848
rect 343048 2836 343054 2848
rect 344554 2836 344560 2848
rect 343048 2808 344560 2836
rect 343048 2796 343054 2808
rect 344554 2796 344560 2808
rect 344612 2796 344618 2848
rect 348050 2796 348056 2848
rect 348108 2836 348114 2848
rect 349154 2836 349160 2848
rect 348108 2808 349160 2836
rect 348108 2796 348114 2808
rect 349154 2796 349160 2808
rect 349212 2796 349218 2848
rect 353938 2796 353944 2848
rect 353996 2836 354002 2848
rect 355226 2836 355232 2848
rect 353996 2808 355232 2836
rect 353996 2796 354002 2808
rect 355226 2796 355232 2808
rect 355284 2796 355290 2848
rect 357434 2796 357440 2848
rect 357492 2836 357498 2848
rect 358722 2836 358728 2848
rect 357492 2808 358728 2836
rect 357492 2796 357498 2808
rect 358722 2796 358728 2808
rect 358780 2796 358786 2848
rect 360838 2796 360844 2848
rect 360896 2836 360902 2848
rect 362310 2836 362316 2848
rect 360896 2808 362316 2836
rect 360896 2796 360902 2808
rect 362310 2796 362316 2808
rect 362368 2796 362374 2848
rect 365806 2796 365812 2848
rect 365864 2836 365870 2848
rect 367094 2836 367100 2848
rect 365864 2808 367100 2836
rect 365864 2796 365870 2808
rect 367094 2796 367100 2808
rect 367152 2796 367158 2848
rect 369394 2796 369400 2848
rect 369452 2836 369458 2848
rect 369854 2836 369860 2848
rect 369452 2808 369860 2836
rect 369452 2796 369458 2808
rect 369854 2796 369860 2808
rect 369912 2796 369918 2848
rect 371878 2796 371884 2848
rect 371936 2836 371942 2848
rect 372890 2836 372896 2848
rect 371936 2808 372896 2836
rect 371936 2796 371942 2808
rect 372890 2796 372896 2808
rect 372948 2796 372954 2848
rect 373994 2796 374000 2848
rect 374052 2836 374058 2848
rect 375282 2836 375288 2848
rect 374052 2808 375288 2836
rect 374052 2796 374058 2808
rect 375282 2796 375288 2808
rect 375340 2796 375346 2848
rect 378778 2796 378784 2848
rect 378836 2836 378842 2848
rect 379974 2836 379980 2848
rect 378836 2808 379980 2836
rect 378836 2796 378842 2808
rect 379974 2796 379980 2808
rect 380032 2796 380038 2848
rect 382274 2796 382280 2848
rect 382332 2836 382338 2848
rect 383562 2836 383568 2848
rect 382332 2808 383568 2836
rect 382332 2796 382338 2808
rect 383562 2796 383568 2808
rect 383620 2796 383626 2848
rect 385678 2796 385684 2848
rect 385736 2836 385742 2848
rect 387150 2836 387156 2848
rect 385736 2808 387156 2836
rect 385736 2796 385742 2808
rect 387150 2796 387156 2808
rect 387208 2796 387214 2848
rect 389818 2796 389824 2848
rect 389876 2836 389882 2848
rect 390646 2836 390652 2848
rect 389876 2808 390652 2836
rect 389876 2796 389882 2808
rect 390646 2796 390652 2808
rect 390704 2796 390710 2848
rect 392670 2796 392676 2848
rect 392728 2836 392734 2848
rect 394234 2836 394240 2848
rect 392728 2808 394240 2836
rect 392728 2796 392734 2808
rect 394234 2796 394240 2808
rect 394292 2796 394298 2848
rect 396644 2836 396672 2876
rect 396718 2864 396724 2916
rect 396776 2904 396782 2916
rect 397730 2904 397736 2916
rect 396776 2876 397736 2904
rect 396776 2864 396782 2876
rect 397730 2864 397736 2876
rect 397788 2864 397794 2916
rect 403618 2864 403624 2916
rect 403676 2904 403682 2916
rect 404814 2904 404820 2916
rect 403676 2876 404820 2904
rect 403676 2864 403682 2876
rect 404814 2864 404820 2876
rect 404872 2864 404878 2916
rect 409340 2904 409368 3012
rect 409432 2972 409460 3080
rect 409509 3043 409567 3049
rect 409509 3009 409521 3043
rect 409555 3040 409567 3043
rect 415486 3040 415492 3052
rect 409555 3012 415492 3040
rect 409555 3009 409567 3012
rect 409509 3003 409567 3009
rect 415486 3000 415492 3012
rect 415544 3000 415550 3052
rect 418126 3040 418154 3080
rect 418798 3068 418804 3120
rect 418856 3108 418862 3120
rect 420178 3108 420184 3120
rect 418856 3080 420184 3108
rect 418856 3068 418862 3080
rect 420178 3068 420184 3080
rect 420236 3068 420242 3120
rect 425440 3108 425468 3216
rect 433242 3204 433248 3216
rect 433300 3204 433306 3256
rect 436738 3204 436744 3256
rect 436796 3204 436802 3256
rect 490558 3204 490564 3256
rect 490616 3244 490622 3256
rect 492306 3244 492312 3256
rect 490616 3216 492312 3244
rect 490616 3204 490622 3216
rect 492306 3204 492312 3216
rect 492364 3204 492370 3256
rect 578602 3204 578608 3256
rect 578660 3244 578666 3256
rect 582929 3247 582987 3253
rect 582929 3244 582941 3247
rect 578660 3216 582941 3244
rect 578660 3204 578666 3216
rect 582929 3213 582941 3216
rect 582975 3213 582987 3247
rect 582929 3207 582987 3213
rect 560938 3136 560944 3188
rect 560996 3176 561002 3188
rect 563238 3176 563244 3188
rect 560996 3148 563244 3176
rect 560996 3136 561002 3148
rect 563238 3136 563244 3148
rect 563296 3136 563302 3188
rect 429654 3108 429660 3120
rect 425440 3080 429660 3108
rect 429654 3068 429660 3080
rect 429712 3068 429718 3120
rect 426158 3040 426164 3052
rect 418126 3012 426164 3040
rect 426158 3000 426164 3012
rect 426216 3000 426222 3052
rect 527818 3000 527824 3052
rect 527876 3040 527882 3052
rect 528646 3040 528652 3052
rect 527876 3012 528652 3040
rect 527876 3000 527882 3012
rect 528646 3000 528652 3012
rect 528704 3000 528710 3052
rect 422570 2972 422576 2984
rect 409432 2944 418154 2972
rect 418126 2904 418154 2944
rect 422266 2944 422576 2972
rect 422266 2904 422294 2944
rect 422570 2932 422576 2944
rect 422628 2932 422634 2984
rect 409340 2876 412036 2904
rect 418126 2876 422294 2904
rect 411898 2836 411904 2848
rect 396644 2808 411904 2836
rect 411898 2796 411904 2808
rect 411956 2796 411962 2848
rect 412008 2836 412036 2876
rect 418982 2836 418988 2848
rect 412008 2808 418988 2836
rect 418982 2796 418988 2808
rect 419040 2796 419046 2848
rect 450078 2796 450084 2848
rect 450136 2836 450142 2848
rect 450906 2836 450912 2848
rect 450136 2808 450912 2836
rect 450136 2796 450142 2808
rect 450906 2796 450912 2808
rect 450964 2796 450970 2848
rect 333882 2768 333888 2780
rect 332612 2740 333888 2768
rect 333882 2728 333888 2740
rect 333940 2728 333946 2780
<< via1 >>
rect 263324 700952 263376 701004
rect 397460 700952 397512 701004
rect 263508 700884 263560 700936
rect 413652 700884 413704 700936
rect 262036 700816 262088 700868
rect 429844 700816 429896 700868
rect 72976 700748 73028 700800
rect 269488 700748 269540 700800
rect 262128 700680 262180 700732
rect 462320 700680 462372 700732
rect 261944 700612 261996 700664
rect 478512 700612 478564 700664
rect 260656 700544 260708 700596
rect 494796 700544 494848 700596
rect 8116 700476 8168 700528
rect 271880 700476 271932 700528
rect 259368 700408 259420 700460
rect 527180 700408 527232 700460
rect 40500 700340 40552 700392
rect 41328 700340 41380 700392
rect 260748 700340 260800 700392
rect 543464 700340 543516 700392
rect 259276 700272 259328 700324
rect 559656 700272 559708 700324
rect 137836 700204 137888 700256
rect 267924 700204 267976 700256
rect 263416 700136 263468 700188
rect 364984 700136 365036 700188
rect 264796 700068 264848 700120
rect 348792 700068 348844 700120
rect 264888 700000 264940 700052
rect 332508 700000 332560 700052
rect 202788 699932 202840 699984
rect 266452 699932 266504 699984
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 170312 699660 170364 699712
rect 171048 699660 171100 699712
rect 235172 699660 235224 699712
rect 235908 699660 235960 699712
rect 266268 699660 266320 699712
rect 267648 699660 267700 699712
rect 257988 696940 258040 696992
rect 580172 696940 580224 696992
rect 259184 683136 259236 683188
rect 580172 683136 580224 683188
rect 257896 670692 257948 670744
rect 580172 670692 580224 670744
rect 3148 656888 3200 656940
rect 273444 656888 273496 656940
rect 256608 643084 256660 643136
rect 580172 643084 580224 643136
rect 257804 630640 257856 630692
rect 580172 630640 580224 630692
rect 256516 616836 256568 616888
rect 580172 616836 580224 616888
rect 3332 605820 3384 605872
rect 274732 605820 274784 605872
rect 255228 590656 255280 590708
rect 579804 590656 579856 590708
rect 255136 576852 255188 576904
rect 580172 576852 580224 576904
rect 255044 563048 255096 563100
rect 579804 563048 579856 563100
rect 3148 553392 3200 553444
rect 276388 553392 276440 553444
rect 253848 536800 253900 536852
rect 580172 536800 580224 536852
rect 253756 524424 253808 524476
rect 580172 524424 580224 524476
rect 252468 510620 252520 510672
rect 580172 510620 580224 510672
rect 3240 500964 3292 501016
rect 277492 500964 277544 501016
rect 252376 484372 252428 484424
rect 580172 484372 580224 484424
rect 252284 470568 252336 470620
rect 579988 470568 580040 470620
rect 251088 456764 251140 456816
rect 580172 456764 580224 456816
rect 3148 448536 3200 448588
rect 278964 448536 279016 448588
rect 250996 430584 251048 430636
rect 580172 430584 580224 430636
rect 250904 418140 250956 418192
rect 580172 418140 580224 418192
rect 249708 404336 249760 404388
rect 580172 404336 580224 404388
rect 2964 397468 3016 397520
rect 281080 397468 281132 397520
rect 3608 380808 3660 380860
rect 274272 380808 274324 380860
rect 3516 380740 3568 380792
rect 273812 380740 273864 380792
rect 3700 380672 3752 380724
rect 275376 380672 275428 380724
rect 3884 380604 3936 380656
rect 276940 380604 276992 380656
rect 3792 380536 3844 380588
rect 276020 380536 276072 380588
rect 3976 380468 4028 380520
rect 277584 380468 277636 380520
rect 4068 380400 4120 380452
rect 278780 380400 278832 380452
rect 3332 380332 3384 380384
rect 279056 380332 279108 380384
rect 3240 380264 3292 380316
rect 280160 380264 280212 380316
rect 3148 380196 3200 380248
rect 280620 380196 280672 380248
rect 3056 380128 3108 380180
rect 281724 380128 281776 380180
rect 41328 380060 41380 380112
rect 271144 380060 271196 380112
rect 106188 379992 106240 380044
rect 269580 379992 269632 380044
rect 89628 379924 89680 379976
rect 270592 379924 270644 379976
rect 154488 379856 154540 379908
rect 269120 379856 269172 379908
rect 171048 379788 171100 379840
rect 219348 379720 219400 379772
rect 258632 379788 258684 379840
rect 259184 379788 259236 379840
rect 260196 379788 260248 379840
rect 260748 379788 260800 379840
rect 261300 379788 261352 379840
rect 262128 379788 262180 379840
rect 262864 379788 262916 379840
rect 263324 379788 263376 379840
rect 250260 379652 250312 379704
rect 250996 379652 251048 379704
rect 251824 379652 251876 379704
rect 252376 379652 252428 379704
rect 253388 379652 253440 379704
rect 253848 379652 253900 379704
rect 254400 379652 254452 379704
rect 255044 379652 255096 379704
rect 256056 379652 256108 379704
rect 256516 379652 256568 379704
rect 257068 379652 257120 379704
rect 257804 379652 257856 379704
rect 267740 379788 267792 379840
rect 268016 379720 268068 379772
rect 280528 379720 280580 379772
rect 290096 379720 290148 379772
rect 264428 379652 264480 379704
rect 264888 379652 264940 379704
rect 265532 379652 265584 379704
rect 299480 379652 299532 379704
rect 235908 379584 235960 379636
rect 254952 379516 255004 379568
rect 255228 379516 255280 379568
rect 263324 379584 263376 379636
rect 263508 379584 263560 379636
rect 266452 379584 266504 379636
rect 271788 379584 271840 379636
rect 283288 379584 283340 379636
rect 266268 379516 266320 379568
rect 282920 379516 282972 379568
rect 234068 379380 234120 379432
rect 283748 379380 283800 379432
rect 243360 379312 243412 379364
rect 295984 379312 296036 379364
rect 232596 379244 232648 379296
rect 285680 379244 285732 379296
rect 231216 379176 231268 379228
rect 287152 379176 287204 379228
rect 248052 379108 248104 379160
rect 302884 379108 302936 379160
rect 222936 379040 222988 379092
rect 284300 379040 284352 379092
rect 242348 378972 242400 379024
rect 304264 378972 304316 379024
rect 228456 378904 228508 378956
rect 291660 378904 291712 378956
rect 245476 378836 245528 378888
rect 307116 378836 307168 378888
rect 246028 378768 246080 378820
rect 314016 378768 314068 378820
rect 249156 378700 249208 378752
rect 318064 378700 318116 378752
rect 215944 378632 215996 378684
rect 287428 378632 287480 378684
rect 213184 378564 213236 378616
rect 292212 378564 292264 378616
rect 3608 378496 3660 378548
rect 282184 378496 282236 378548
rect 248236 378428 248288 378480
rect 580172 378428 580224 378480
rect 239680 378360 239732 378412
rect 240048 378292 240100 378344
rect 237196 378224 237248 378276
rect 237104 378156 237156 378208
rect 244924 377884 244976 377936
rect 246580 377816 246632 377868
rect 300216 377816 300268 377868
rect 243912 377748 243964 377800
rect 298836 377748 298888 377800
rect 224224 377680 224276 377732
rect 282920 377680 282972 377732
rect 246948 377612 247000 377664
rect 238576 377587 238628 377596
rect 238576 377553 238585 377587
rect 238585 377553 238619 377587
rect 238619 377553 238628 377587
rect 238576 377544 238628 377553
rect 239220 377587 239272 377596
rect 239220 377553 239229 377587
rect 239229 377553 239263 377587
rect 239263 377553 239272 377587
rect 239220 377544 239272 377553
rect 240784 377587 240836 377596
rect 240784 377553 240793 377587
rect 240793 377553 240827 377587
rect 240827 377553 240836 377587
rect 240784 377544 240836 377553
rect 241612 377587 241664 377596
rect 241612 377553 241621 377587
rect 241621 377553 241655 377587
rect 241655 377553 241664 377587
rect 241612 377544 241664 377553
rect 247592 377587 247644 377596
rect 247592 377553 247601 377587
rect 247601 377553 247635 377587
rect 247635 377553 247644 377587
rect 247592 377544 247644 377553
rect 305644 377612 305696 377664
rect 309784 377544 309836 377596
rect 3516 377476 3568 377528
rect 271788 377476 271840 377528
rect 3424 377408 3476 377460
rect 280528 377408 280580 377460
rect 284852 377451 284904 377460
rect 284852 377417 284861 377451
rect 284861 377417 284895 377451
rect 284895 377417 284904 377451
rect 284852 377408 284904 377417
rect 220176 377340 220228 377392
rect 285864 377340 285916 377392
rect 288532 377383 288584 377392
rect 288532 377349 288541 377383
rect 288541 377349 288575 377383
rect 288575 377349 288584 377383
rect 288532 377340 288584 377349
rect 290648 377383 290700 377392
rect 290648 377349 290657 377383
rect 290657 377349 290691 377383
rect 290691 377349 290700 377383
rect 290648 377340 290700 377349
rect 293224 377340 293276 377392
rect 226984 377272 227036 377324
rect 316684 377204 316736 377256
rect 214564 377136 214616 377188
rect 209044 377068 209096 377120
rect 4804 377000 4856 377052
rect 318064 365644 318116 365696
rect 580172 365644 580224 365696
rect 302884 353200 302936 353252
rect 580172 353200 580224 353252
rect 3148 346332 3200 346384
rect 224224 346332 224276 346384
rect 125508 337628 125560 337680
rect 238990 337900 239042 337952
rect 239358 337900 239410 337952
rect 234804 337832 234856 337884
rect 235586 337832 235638 337884
rect 238622 337832 238674 337884
rect 237932 337628 237984 337680
rect 239036 337764 239088 337816
rect 239220 337628 239272 337680
rect 242026 337832 242078 337884
rect 243222 337832 243274 337884
rect 243360 337832 243412 337884
rect 241520 337628 241572 337680
rect 242900 337628 242952 337680
rect 243084 337628 243136 337680
rect 122104 337560 122156 337612
rect 97908 337492 97960 337544
rect 244970 337900 245022 337952
rect 246074 337900 246126 337952
rect 246626 337900 246678 337952
rect 247270 337900 247322 337952
rect 247730 337900 247782 337952
rect 251134 337900 251186 337952
rect 262956 337900 263008 337952
rect 263830 337900 263882 337952
rect 264198 337900 264250 337952
rect 264566 337900 264618 337952
rect 274410 337900 274462 337952
rect 276342 337900 276394 337952
rect 276710 337900 276762 337952
rect 277078 337900 277130 337952
rect 281218 337900 281270 337952
rect 283656 337943 283708 337952
rect 283656 337909 283665 337943
rect 283665 337909 283699 337943
rect 283699 337909 283708 337943
rect 283656 337900 283708 337909
rect 283978 337900 284030 337952
rect 290602 337900 290654 337952
rect 294466 337900 294518 337952
rect 294972 337900 295024 337952
rect 245062 337764 245114 337816
rect 246166 337832 246218 337884
rect 245752 337628 245804 337680
rect 246028 337628 246080 337680
rect 247316 337764 247368 337816
rect 248098 337764 248150 337816
rect 250904 337764 250956 337816
rect 247132 337628 247184 337680
rect 250720 337628 250772 337680
rect 250904 337628 250956 337680
rect 251502 337832 251554 337884
rect 251778 337832 251830 337884
rect 251732 337628 251784 337680
rect 253112 337832 253164 337884
rect 253618 337832 253670 337884
rect 253710 337832 253762 337884
rect 256010 337832 256062 337884
rect 253112 337696 253164 337748
rect 253388 337628 253440 337680
rect 253572 337628 253624 337680
rect 255642 337764 255694 337816
rect 255688 337628 255740 337680
rect 261254 337832 261306 337884
rect 258678 337764 258730 337816
rect 260840 337764 260892 337816
rect 257436 337628 257488 337680
rect 264796 337832 264848 337884
rect 269902 337832 269954 337884
rect 270638 337832 270690 337884
rect 271466 337832 271518 337884
rect 272570 337832 272622 337884
rect 278182 337832 278234 337884
rect 280022 337832 280074 337884
rect 293638 337832 293690 337884
rect 294650 337832 294702 337884
rect 294880 337832 294932 337884
rect 263048 337628 263100 337680
rect 264704 337628 264756 337680
rect 280942 337764 280994 337816
rect 281172 337764 281224 337816
rect 284346 337764 284398 337816
rect 285082 337764 285134 337816
rect 286186 337764 286238 337816
rect 270776 337628 270828 337680
rect 349160 337628 349212 337680
rect 272248 337560 272300 337612
rect 360844 337560 360896 337612
rect 273444 337535 273496 337544
rect 273444 337501 273453 337535
rect 273453 337501 273487 337535
rect 273487 337501 273496 337535
rect 273444 337492 273496 337501
rect 367100 337492 367152 337544
rect 91008 337424 91060 337476
rect 244188 337424 244240 337476
rect 272892 337424 272944 337476
rect 369860 337424 369912 337476
rect 86868 337356 86920 337408
rect 243820 337356 243872 337408
rect 278964 337356 279016 337408
rect 425704 337356 425756 337408
rect 81348 337288 81400 337340
rect 242900 337288 242952 337340
rect 279056 337288 279108 337340
rect 427820 337288 427872 337340
rect 70308 337220 70360 337272
rect 241520 337220 241572 337272
rect 279424 337220 279476 337272
rect 432052 337220 432104 337272
rect 66168 337152 66220 337204
rect 241704 337152 241756 337204
rect 280436 337195 280488 337204
rect 280436 337161 280445 337195
rect 280445 337161 280479 337195
rect 280479 337161 280488 337195
rect 280436 337152 280488 337161
rect 436744 337152 436796 337204
rect 50344 337084 50396 337136
rect 239496 337084 239548 337136
rect 283288 337084 283340 337136
rect 468484 337084 468536 337136
rect 48228 337016 48280 337068
rect 239864 337016 239916 337068
rect 283472 337016 283524 337068
rect 470600 337016 470652 337068
rect 41328 336948 41380 337000
rect 239128 336948 239180 337000
rect 472624 336948 472676 337000
rect 34428 336880 34480 336932
rect 238392 336880 238444 336932
rect 292948 336880 293000 336932
rect 560944 336880 560996 336932
rect 29644 336812 29696 336864
rect 237656 336812 237708 336864
rect 294144 336812 294196 336864
rect 574100 336812 574152 336864
rect 12348 336744 12400 336796
rect 236184 336744 236236 336796
rect 224224 336676 224276 336728
rect 251916 336676 251968 336728
rect 253572 336676 253624 336728
rect 263416 336676 263468 336728
rect 280712 336744 280764 336796
rect 280896 336744 280948 336796
rect 284852 336744 284904 336796
rect 285036 336744 285088 336796
rect 294972 336744 295024 336796
rect 260656 336608 260708 336660
rect 262312 336608 262364 336660
rect 262496 336608 262548 336660
rect 233056 336540 233108 336592
rect 261024 336540 261076 336592
rect 228364 336472 228416 336524
rect 258080 336472 258132 336524
rect 262496 336472 262548 336524
rect 263600 336472 263652 336524
rect 222844 336404 222896 336456
rect 206284 336336 206336 336388
rect 252560 336404 252612 336456
rect 252652 336404 252704 336456
rect 256148 336404 256200 336456
rect 262220 336404 262272 336456
rect 263876 336404 263928 336456
rect 256976 336336 257028 336388
rect 264704 336676 264756 336728
rect 298744 336676 298796 336728
rect 272616 336608 272668 336660
rect 273168 336608 273220 336660
rect 285864 336608 285916 336660
rect 320824 336608 320876 336660
rect 266544 336540 266596 336592
rect 285128 336540 285180 336592
rect 286968 336540 287020 336592
rect 322204 336540 322256 336592
rect 265808 336472 265860 336524
rect 286600 336472 286652 336524
rect 287336 336472 287388 336524
rect 323676 336472 323728 336524
rect 265440 336404 265492 336456
rect 282644 336404 282696 336456
rect 282828 336404 282880 336456
rect 289084 336404 289136 336456
rect 331864 336404 331916 336456
rect 277492 336336 277544 336388
rect 204904 336268 204956 336320
rect 266912 336268 266964 336320
rect 273812 336268 273864 336320
rect 274364 336268 274416 336320
rect 277400 336268 277452 336320
rect 323584 336336 323636 336388
rect 336004 336268 336056 336320
rect 198004 336200 198056 336252
rect 202144 336132 202196 336184
rect 196624 336064 196676 336116
rect 252560 336200 252612 336252
rect 258816 336200 258868 336252
rect 265164 336200 265216 336252
rect 376024 336200 376076 336252
rect 251272 336132 251324 336184
rect 251456 336132 251508 336184
rect 251824 336132 251876 336184
rect 260012 336132 260064 336184
rect 268660 336132 268712 336184
rect 393964 336132 394016 336184
rect 254032 336064 254084 336116
rect 263048 336064 263100 336116
rect 284300 336064 284352 336116
rect 285956 336064 286008 336116
rect 497464 336064 497516 336116
rect 195244 335996 195296 336048
rect 253020 335996 253072 336048
rect 265256 335996 265308 336048
rect 272892 335996 272944 336048
rect 231768 335928 231820 335980
rect 260380 335928 260432 335980
rect 266084 335928 266136 335980
rect 231124 335860 231176 335912
rect 254768 335860 254820 335912
rect 262956 335860 263008 335912
rect 267004 335860 267056 335912
rect 232504 335792 232556 335844
rect 255136 335792 255188 335844
rect 272892 335792 272944 335844
rect 233976 335724 234028 335776
rect 258448 335724 258500 335776
rect 286968 335996 287020 336048
rect 287704 335996 287756 336048
rect 294972 335996 295024 336048
rect 295248 335996 295300 336048
rect 522304 335996 522356 336048
rect 289544 335928 289596 335980
rect 303252 335928 303304 335980
rect 294604 335860 294656 335912
rect 295156 335860 295208 335912
rect 295708 335860 295760 335912
rect 282828 335792 282880 335844
rect 287520 335792 287572 335844
rect 288072 335792 288124 335844
rect 299480 335792 299532 335844
rect 276940 335724 276992 335776
rect 278320 335724 278372 335776
rect 285220 335724 285272 335776
rect 285496 335767 285548 335776
rect 285496 335733 285505 335767
rect 285505 335733 285539 335767
rect 285539 335733 285548 335767
rect 285496 335724 285548 335733
rect 286508 335724 286560 335776
rect 296628 335724 296680 335776
rect 233884 335656 233936 335708
rect 234436 335588 234488 335640
rect 259184 335656 259236 335708
rect 269580 335656 269632 335708
rect 254400 335588 254452 335640
rect 266728 335588 266780 335640
rect 278504 335656 278556 335708
rect 278688 335656 278740 335708
rect 279516 335656 279568 335708
rect 279700 335656 279752 335708
rect 230480 335520 230532 335572
rect 252284 335520 252336 335572
rect 253848 335520 253900 335572
rect 262312 335520 262364 335572
rect 268016 335520 268068 335572
rect 278320 335520 278372 335572
rect 233148 335452 233200 335504
rect 233424 335384 233476 335436
rect 257344 335452 257396 335504
rect 260104 335452 260156 335504
rect 261300 335452 261352 335504
rect 262772 335452 262824 335504
rect 263508 335452 263560 335504
rect 269764 335452 269816 335504
rect 270132 335452 270184 335504
rect 271972 335452 272024 335504
rect 272892 335452 272944 335504
rect 273352 335452 273404 335504
rect 231676 335316 231728 335368
rect 253296 335384 253348 335436
rect 257712 335384 257764 335436
rect 260656 335384 260708 335436
rect 261760 335384 261812 335436
rect 262588 335384 262640 335436
rect 263416 335384 263468 335436
rect 265072 335384 265124 335436
rect 265808 335384 265860 335436
rect 268660 335384 268712 335436
rect 269028 335384 269080 335436
rect 271328 335384 271380 335436
rect 271696 335384 271748 335436
rect 272340 335384 272392 335436
rect 273076 335384 273128 335436
rect 254860 335316 254912 335368
rect 255780 335316 255832 335368
rect 258724 335316 258776 335368
rect 259736 335316 259788 335368
rect 261116 335316 261168 335368
rect 261852 335316 261904 335368
rect 266636 335316 266688 335368
rect 267096 335316 267148 335368
rect 267280 335316 267332 335368
rect 267832 335316 267884 335368
rect 268200 335316 268252 335368
rect 151728 335248 151780 335300
rect 250444 335248 250496 335300
rect 147588 335180 147640 335232
rect 250076 335180 250128 335232
rect 262128 335180 262180 335232
rect 262864 335180 262916 335232
rect 268752 335316 268804 335368
rect 268936 335316 268988 335368
rect 270500 335316 270552 335368
rect 270960 335316 271012 335368
rect 271236 335316 271288 335368
rect 271512 335316 271564 335368
rect 271880 335316 271932 335368
rect 273628 335316 273680 335368
rect 274088 335316 274140 335368
rect 277676 335452 277728 335504
rect 278504 335452 278556 335504
rect 275192 335384 275244 335436
rect 274640 335316 274692 335368
rect 275468 335316 275520 335368
rect 275928 335316 275980 335368
rect 271696 335248 271748 335300
rect 274456 335248 274508 335300
rect 268752 335180 268804 335232
rect 276756 335384 276808 335436
rect 277308 335384 277360 335436
rect 278136 335316 278188 335368
rect 278412 335316 278464 335368
rect 279148 335384 279200 335436
rect 279884 335384 279936 335436
rect 280804 335384 280856 335436
rect 281448 335384 281500 335436
rect 278780 335316 278832 335368
rect 279516 335316 279568 335368
rect 282184 335316 282236 335368
rect 282460 335316 282512 335368
rect 288808 335656 288860 335708
rect 292764 335656 292816 335708
rect 304172 335792 304224 335844
rect 282828 335588 282880 335640
rect 285496 335520 285548 335572
rect 287244 335520 287296 335572
rect 287980 335520 288032 335572
rect 284392 335452 284444 335504
rect 284484 335452 284536 335504
rect 285404 335452 285456 335504
rect 287612 335452 287664 335504
rect 288072 335452 288124 335504
rect 285680 335384 285732 335436
rect 286324 335427 286376 335436
rect 286324 335393 286333 335427
rect 286333 335393 286367 335427
rect 286367 335393 286376 335427
rect 286324 335384 286376 335393
rect 287244 335384 287296 335436
rect 287888 335384 287940 335436
rect 284668 335316 284720 335368
rect 285404 335316 285456 335368
rect 285772 335316 285824 335368
rect 286876 335316 286928 335368
rect 287704 335316 287756 335368
rect 288256 335316 288308 335368
rect 289176 335588 289228 335640
rect 296536 335588 296588 335640
rect 294880 335520 294932 335572
rect 295248 335520 295300 335572
rect 298192 335520 298244 335572
rect 288624 335452 288676 335504
rect 289452 335452 289504 335504
rect 289912 335452 289964 335504
rect 288992 335384 289044 335436
rect 289544 335384 289596 335436
rect 294236 335384 294288 335436
rect 294880 335384 294932 335436
rect 295432 335384 295484 335436
rect 288900 335316 288952 335368
rect 289360 335316 289412 335368
rect 290096 335316 290148 335368
rect 290924 335316 290976 335368
rect 291752 335316 291804 335368
rect 292120 335316 292172 335368
rect 292580 335316 292632 335368
rect 292672 335316 292724 335368
rect 293868 335316 293920 335368
rect 294788 335316 294840 335368
rect 295156 335316 295208 335368
rect 296352 335316 296404 335368
rect 387800 335248 387852 335300
rect 394700 335180 394752 335232
rect 144828 335112 144880 335164
rect 249708 335112 249760 335164
rect 277768 335112 277820 335164
rect 414664 335112 414716 335164
rect 126888 335044 126940 335096
rect 234528 335044 234580 335096
rect 140688 334976 140740 335028
rect 249340 335044 249392 335096
rect 279608 335044 279660 335096
rect 432604 335044 432656 335096
rect 263968 334976 264020 335028
rect 264796 334976 264848 335028
rect 284760 334976 284812 335028
rect 137284 334908 137336 334960
rect 248972 334908 249024 334960
rect 480260 334976 480312 335028
rect 483020 334908 483072 334960
rect 133788 334840 133840 334892
rect 248604 334840 248656 334892
rect 487160 334840 487212 334892
rect 129004 334772 129056 334824
rect 247960 334772 248012 334824
rect 287520 334772 287572 334824
rect 296628 334772 296680 334824
rect 500960 334772 501012 334824
rect 87604 334704 87656 334756
rect 243636 334704 243688 334756
rect 257344 334704 257396 334756
rect 260012 334704 260064 334756
rect 282092 334704 282144 334756
rect 282368 334704 282420 334756
rect 284392 334704 284444 334756
rect 299388 334704 299440 334756
rect 299480 334704 299532 334756
rect 514760 334704 514812 334756
rect 52368 334636 52420 334688
rect 240232 334636 240284 334688
rect 273260 334636 273312 334688
rect 17868 334568 17920 334620
rect 236644 334568 236696 334620
rect 237472 334568 237524 334620
rect 237748 334568 237800 334620
rect 239128 334568 239180 334620
rect 239680 334568 239732 334620
rect 242992 334568 243044 334620
rect 243452 334568 243504 334620
rect 244924 334568 244976 334620
rect 245200 334568 245252 334620
rect 246396 334568 246448 334620
rect 246580 334568 246632 334620
rect 251640 334568 251692 334620
rect 252468 334568 252520 334620
rect 252836 334568 252888 334620
rect 253756 334568 253808 334620
rect 258356 334568 258408 334620
rect 259368 334568 259420 334620
rect 260012 334568 260064 334620
rect 260748 334568 260800 334620
rect 273628 334568 273680 334620
rect 273996 334568 274048 334620
rect 282092 334568 282144 334620
rect 282736 334568 282788 334620
rect 155224 334500 155276 334552
rect 250812 334500 250864 334552
rect 271328 334543 271380 334552
rect 271328 334509 271337 334543
rect 271337 334509 271371 334543
rect 271371 334509 271380 334543
rect 271328 334500 271380 334509
rect 275560 334500 275612 334552
rect 275836 334500 275888 334552
rect 285496 334636 285548 334688
rect 295340 334636 295392 334688
rect 296536 334636 296588 334688
rect 532700 334636 532752 334688
rect 290004 334568 290056 334620
rect 535460 334568 535512 334620
rect 371884 334500 371936 334552
rect 158628 334432 158680 334484
rect 250904 334432 250956 334484
rect 271052 334432 271104 334484
rect 351920 334432 351972 334484
rect 161388 334364 161440 334416
rect 233148 334364 233200 334416
rect 169668 334296 169720 334348
rect 230480 334296 230532 334348
rect 233240 334296 233292 334348
rect 252560 334364 252612 334416
rect 262404 334364 262456 334416
rect 263416 334364 263468 334416
rect 263784 334364 263836 334416
rect 264244 334364 264296 334416
rect 269212 334364 269264 334416
rect 333980 334364 334032 334416
rect 268384 334296 268436 334348
rect 324320 334296 324372 334348
rect 194416 334228 194468 334280
rect 254768 334228 254820 334280
rect 267556 334228 267608 334280
rect 316040 334228 316092 334280
rect 212448 334160 212500 334212
rect 256792 334160 256844 334212
rect 267188 334160 267240 334212
rect 313280 334160 313332 334212
rect 220084 334092 220136 334144
rect 257528 334092 257580 334144
rect 286600 334092 286652 334144
rect 309140 334092 309192 334144
rect 227628 334024 227680 334076
rect 258264 334024 258316 334076
rect 285128 334024 285180 334076
rect 306380 334024 306432 334076
rect 230388 333956 230440 334008
rect 258540 333956 258592 334008
rect 286968 333956 287020 334008
rect 302240 333956 302292 334008
rect 187608 333888 187660 333940
rect 254216 333888 254268 333940
rect 418804 333888 418856 333940
rect 166908 333820 166960 333872
rect 252008 333820 252060 333872
rect 278688 333820 278740 333872
rect 423680 333820 423732 333872
rect 162768 333752 162820 333804
rect 251916 333752 251968 333804
rect 287336 333752 287388 333804
rect 465172 333752 465224 333804
rect 144736 333684 144788 333736
rect 249800 333684 249852 333736
rect 292120 333684 292172 333736
rect 292488 333684 292540 333736
rect 292580 333684 292632 333736
rect 489920 333684 489972 333736
rect 135168 333616 135220 333668
rect 248696 333616 248748 333668
rect 265624 333616 265676 333668
rect 298100 333616 298152 333668
rect 298192 333616 298244 333668
rect 507860 333616 507912 333668
rect 88984 333548 89036 333600
rect 244004 333548 244056 333600
rect 287060 333548 287112 333600
rect 506480 333548 506532 333600
rect 83464 333480 83516 333532
rect 239312 333480 239364 333532
rect 265992 333480 266044 333532
rect 300124 333480 300176 333532
rect 303252 333480 303304 333532
rect 529940 333480 529992 333532
rect 73068 333412 73120 333464
rect 242440 333412 242492 333464
rect 288808 333412 288860 333464
rect 524512 333412 524564 333464
rect 59268 333344 59320 333396
rect 240968 333344 241020 333396
rect 290740 333344 290792 333396
rect 542452 333344 542504 333396
rect 55128 333276 55180 333328
rect 240600 333276 240652 333328
rect 280620 333276 280672 333328
rect 281264 333276 281316 333328
rect 283196 333276 283248 333328
rect 283748 333276 283800 333328
rect 291200 333276 291252 333328
rect 292304 333276 292356 333328
rect 296444 333276 296496 333328
rect 547880 333276 547932 333328
rect 22008 333208 22060 333260
rect 237196 333208 237248 333260
rect 258816 333208 258868 333260
rect 259828 333208 259880 333260
rect 264060 333208 264112 333260
rect 264520 333208 264572 333260
rect 265532 333208 265584 333260
rect 266084 333208 266136 333260
rect 272708 333208 272760 333260
rect 273168 333208 273220 333260
rect 273904 333208 273956 333260
rect 274180 333208 274232 333260
rect 276480 333208 276532 333260
rect 277124 333208 277176 333260
rect 277584 333208 277636 333260
rect 278320 333208 278372 333260
rect 280252 333208 280304 333260
rect 281448 333208 281500 333260
rect 283564 333208 283616 333260
rect 284024 333208 284076 333260
rect 298008 333208 298060 333260
rect 568580 333208 568632 333260
rect 169576 333140 169628 333192
rect 252376 333140 252428 333192
rect 405740 333140 405792 333192
rect 191748 333072 191800 333124
rect 254584 333072 254636 333124
rect 412640 333072 412692 333124
rect 198648 333004 198700 333056
rect 255228 333004 255280 333056
rect 285220 333004 285272 333056
rect 398840 333004 398892 333056
rect 179328 332936 179380 332988
rect 233424 332936 233476 332988
rect 254584 332936 254636 332988
rect 259092 332936 259144 332988
rect 353944 332936 353996 332988
rect 206928 332868 206980 332920
rect 252652 332868 252704 332920
rect 269304 332868 269356 332920
rect 331956 332868 332008 332920
rect 210976 332800 211028 332852
rect 256516 332800 256568 332852
rect 268108 332800 268160 332852
rect 321560 332800 321612 332852
rect 216588 332732 216640 332784
rect 257160 332732 257212 332784
rect 266912 332732 266964 332784
rect 310520 332732 310572 332784
rect 223488 332664 223540 332716
rect 257804 332664 257856 332716
rect 266728 332664 266780 332716
rect 307024 332664 307076 332716
rect 227536 332596 227588 332648
rect 258172 332596 258224 332648
rect 153108 332528 153160 332580
rect 250536 332528 250588 332580
rect 284852 332528 284904 332580
rect 430580 332528 430632 332580
rect 148968 332460 149020 332512
rect 250168 332460 250220 332512
rect 476120 332460 476172 332512
rect 142068 332392 142120 332444
rect 249432 332392 249484 332444
rect 284576 332392 284628 332444
rect 481640 332392 481692 332444
rect 137928 332324 137980 332376
rect 249064 332324 249116 332376
rect 285036 332324 285088 332376
rect 484400 332324 484452 332376
rect 124128 332256 124180 332308
rect 247592 332256 247644 332308
rect 286232 332256 286284 332308
rect 499672 332256 499724 332308
rect 104808 332188 104860 332240
rect 245660 332188 245712 332240
rect 287428 332188 287480 332240
rect 510712 332188 510764 332240
rect 95148 332120 95200 332172
rect 244648 332120 244700 332172
rect 296352 332120 296404 332172
rect 525800 332120 525852 332172
rect 77208 332052 77260 332104
rect 62028 331984 62080 332036
rect 241336 332052 241388 332104
rect 288532 332052 288584 332104
rect 520280 332052 520332 332104
rect 53104 331916 53156 331968
rect 239956 331984 240008 332036
rect 539692 331984 539744 332036
rect 32404 331848 32456 331900
rect 238024 331916 238076 331968
rect 290372 331916 290424 331968
rect 538220 331916 538272 331968
rect 287060 331848 287112 331900
rect 295524 331848 295576 331900
rect 547972 331848 548024 331900
rect 155868 331780 155920 331832
rect 250720 331780 250772 331832
rect 274824 331780 274876 331832
rect 385684 331780 385736 331832
rect 184848 331712 184900 331764
rect 253940 331712 253992 331764
rect 271696 331712 271748 331764
rect 357440 331712 357492 331764
rect 188988 331644 189040 331696
rect 254308 331644 254360 331696
rect 269672 331644 269724 331696
rect 338120 331644 338172 331696
rect 213828 331576 213880 331628
rect 256884 331576 256936 331628
rect 276940 331576 276992 331628
rect 335360 331576 335412 331628
rect 224868 331508 224920 331560
rect 257988 331508 258040 331560
rect 268476 331508 268528 331560
rect 324412 331508 324464 331560
rect 234344 331440 234396 331492
rect 258908 331440 258960 331492
rect 267372 331440 267424 331492
rect 313924 331440 313976 331492
rect 242716 331372 242768 331424
rect 266360 331372 266412 331424
rect 305000 331372 305052 331424
rect 193128 331168 193180 331220
rect 254676 331168 254728 331220
rect 279792 331168 279844 331220
rect 434720 331168 434772 331220
rect 153016 331100 153068 331152
rect 250628 331100 250680 331152
rect 293040 331100 293092 331152
rect 450544 331100 450596 331152
rect 111708 331032 111760 331084
rect 246580 331032 246632 331084
rect 285312 331032 285364 331084
rect 488540 331032 488592 331084
rect 108948 330964 109000 331016
rect 245752 330964 245804 331016
rect 102048 330896 102100 330948
rect 245292 330896 245344 330948
rect 79324 330828 79376 330880
rect 242808 330828 242860 330880
rect 284300 330964 284352 331016
rect 285588 330964 285640 331016
rect 490564 330964 490616 331016
rect 286692 330896 286744 330948
rect 502340 330896 502392 330948
rect 287796 330828 287848 330880
rect 512644 330828 512696 330880
rect 68284 330760 68336 330812
rect 241796 330760 241848 330812
rect 272892 330760 272944 330812
rect 299940 330760 299992 330812
rect 536840 330760 536892 330812
rect 57244 330692 57296 330744
rect 240324 330692 240376 330744
rect 39304 330624 39356 330676
rect 238944 330624 238996 330676
rect 37188 330556 37240 330608
rect 22744 330488 22796 330540
rect 236276 330556 236328 330608
rect 255596 330488 255648 330540
rect 256240 330488 256292 330540
rect 258632 330488 258684 330540
rect 259276 330488 259328 330540
rect 267188 330488 267240 330540
rect 267464 330488 267516 330540
rect 195888 330420 195940 330472
rect 255044 330420 255096 330472
rect 255412 330420 255464 330472
rect 255964 330420 256016 330472
rect 259644 330420 259696 330472
rect 260288 330420 260340 330472
rect 272156 330420 272208 330472
rect 272800 330420 272852 330472
rect 289268 330692 289320 330744
rect 528652 330692 528704 330744
rect 291108 330624 291160 330676
rect 546500 330624 546552 330676
rect 293316 330556 293368 330608
rect 294052 330488 294104 330540
rect 294788 330488 294840 330540
rect 295800 330556 295852 330608
rect 564532 330556 564584 330608
rect 565820 330488 565872 330540
rect 273076 330420 273128 330472
rect 274088 330420 274140 330472
rect 375380 330420 375432 330472
rect 202788 330352 202840 330404
rect 254860 330352 254912 330404
rect 217968 330284 218020 330336
rect 257252 330352 257304 330404
rect 270408 330352 270460 330404
rect 342904 330352 342956 330404
rect 255780 330327 255832 330336
rect 255780 330293 255789 330327
rect 255789 330293 255823 330327
rect 255823 330293 255832 330327
rect 255780 330284 255832 330293
rect 255872 330284 255924 330336
rect 256332 330284 256384 330336
rect 260840 330284 260892 330336
rect 261116 330284 261168 330336
rect 268936 330284 268988 330336
rect 328460 330284 328512 330336
rect 220728 330216 220780 330268
rect 238576 330148 238628 330200
rect 255412 330216 255464 330268
rect 256608 330216 256660 330268
rect 267648 330216 267700 330268
rect 317420 330216 317472 330268
rect 257620 330148 257672 330200
rect 261116 330148 261168 330200
rect 261576 330148 261628 330200
rect 263876 330148 263928 330200
rect 264244 330148 264296 330200
rect 275100 329740 275152 329792
rect 389824 329740 389876 329792
rect 146208 329672 146260 329724
rect 249984 329672 250036 329724
rect 276848 329672 276900 329724
rect 407120 329672 407172 329724
rect 99288 329604 99340 329656
rect 277216 329604 277268 329656
rect 409880 329604 409932 329656
rect 93124 329536 93176 329588
rect 244372 329536 244424 329588
rect 280068 329536 280120 329588
rect 438860 329536 438912 329588
rect 75184 329468 75236 329520
rect 242532 329468 242584 329520
rect 283656 329468 283708 329520
rect 474740 329468 474792 329520
rect 71044 329400 71096 329452
rect 242164 329400 242216 329452
rect 288256 329400 288308 329452
rect 517520 329400 517572 329452
rect 63408 329332 63460 329384
rect 241428 329332 241480 329384
rect 289636 329332 289688 329384
rect 530584 329332 530636 329384
rect 61384 329264 61436 329316
rect 241060 329264 241112 329316
rect 304172 329264 304224 329316
rect 561680 329264 561732 329316
rect 57336 329196 57388 329248
rect 240692 329196 240744 329248
rect 291844 329196 291896 329248
rect 551284 329196 551336 329248
rect 39396 329128 39448 329180
rect 236828 329128 236880 329180
rect 291752 329128 291804 329180
rect 556160 329128 556212 329180
rect 32496 329060 32548 329112
rect 238116 329060 238168 329112
rect 264888 329060 264940 329112
rect 291200 329060 291252 329112
rect 569960 329060 570012 329112
rect 273628 328992 273680 329044
rect 378784 328992 378836 329044
rect 270040 328924 270092 328976
rect 340880 328924 340932 328976
rect 270132 328695 270184 328704
rect 270132 328661 270141 328695
rect 270141 328661 270175 328695
rect 270175 328661 270184 328695
rect 270132 328652 270184 328661
rect 273444 328380 273496 328432
rect 382280 328380 382332 328432
rect 275744 328312 275796 328364
rect 392584 328312 392636 328364
rect 265900 328244 265952 328296
rect 266176 328244 266228 328296
rect 278320 328244 278372 328296
rect 414020 328244 414072 328296
rect 119988 328176 120040 328228
rect 245108 328176 245160 328228
rect 277860 328176 277912 328228
rect 416780 328176 416832 328228
rect 113088 328108 113140 328160
rect 246396 328108 246448 328160
rect 278228 328108 278280 328160
rect 420920 328108 420972 328160
rect 111064 328040 111116 328092
rect 246028 328040 246080 328092
rect 293684 328040 293736 328092
rect 453304 328040 453356 328092
rect 106188 327972 106240 328024
rect 245844 327972 245896 328024
rect 290924 327972 290976 328024
rect 464344 327972 464396 328024
rect 95056 327904 95108 327956
rect 244740 327904 244792 327956
rect 286508 327904 286560 327956
rect 466460 327904 466512 327956
rect 43444 327836 43496 327888
rect 237288 327836 237340 327888
rect 284116 327836 284168 327888
rect 477500 327836 477552 327888
rect 45468 327768 45520 327820
rect 239312 327768 239364 327820
rect 286784 327768 286836 327820
rect 503720 327768 503772 327820
rect 28908 327700 28960 327752
rect 237472 327700 237524 327752
rect 292120 327700 292172 327752
rect 560300 327700 560352 327752
rect 275560 326884 275612 326936
rect 396724 326884 396776 326936
rect 278596 326816 278648 326868
rect 423772 326816 423824 326868
rect 285404 326748 285456 326800
rect 293592 326748 293644 326800
rect 443644 326748 443696 326800
rect 234988 326723 235040 326732
rect 234988 326689 234997 326723
rect 234997 326689 235031 326723
rect 235031 326689 235040 326723
rect 234988 326680 235040 326689
rect 241612 326680 241664 326732
rect 284944 326680 284996 326732
rect 117228 326612 117280 326664
rect 246856 326612 246908 326664
rect 68376 326544 68428 326596
rect 58624 326476 58676 326528
rect 240876 326544 240928 326596
rect 280620 326587 280672 326596
rect 280620 326553 280629 326587
rect 280629 326553 280663 326587
rect 280663 326553 280672 326587
rect 280620 326544 280672 326553
rect 286876 326544 286928 326596
rect 290556 326680 290608 326732
rect 461584 326680 461636 326732
rect 481732 326612 481784 326664
rect 50988 326408 51040 326460
rect 240048 326476 240100 326528
rect 288072 326476 288124 326528
rect 485780 326544 485832 326596
rect 35808 326340 35860 326392
rect 238484 326408 238536 326460
rect 243084 326408 243136 326460
rect 244096 326408 244148 326460
rect 273812 326408 273864 326460
rect 274548 326408 274600 326460
rect 281356 326408 281408 326460
rect 282368 326408 282420 326460
rect 282552 326408 282604 326460
rect 289452 326408 289504 326460
rect 492680 326476 492732 326528
rect 236184 326340 236236 326392
rect 236552 326340 236604 326392
rect 237380 326340 237432 326392
rect 237932 326340 237984 326392
rect 239036 326340 239088 326392
rect 239404 326340 239456 326392
rect 243176 326340 243228 326392
rect 243728 326340 243780 326392
rect 246120 326340 246172 326392
rect 246948 326340 247000 326392
rect 247132 326340 247184 326392
rect 248236 326340 248288 326392
rect 248696 326340 248748 326392
rect 249156 326340 249208 326392
rect 273536 326340 273588 326392
rect 273996 326340 274048 326392
rect 275008 326340 275060 326392
rect 275376 326340 275428 326392
rect 280344 326340 280396 326392
rect 280988 326340 281040 326392
rect 280620 326315 280672 326324
rect 280620 326281 280629 326315
rect 280629 326281 280663 326315
rect 280663 326281 280672 326315
rect 280620 326272 280672 326281
rect 235172 326204 235224 326256
rect 235632 326204 235684 326256
rect 247224 326204 247276 326256
rect 247408 326204 247460 326256
rect 247500 326204 247552 326256
rect 247684 326204 247736 326256
rect 288992 326340 289044 326392
rect 289728 326340 289780 326392
rect 506572 326408 506624 326460
rect 519544 326340 519596 326392
rect 281448 326204 281500 326256
rect 282276 326204 282328 326256
rect 282644 326204 282696 326256
rect 281724 326136 281776 326188
rect 282828 326136 282880 326188
rect 247224 326068 247276 326120
rect 248328 326068 248380 326120
rect 281816 326068 281868 326120
rect 282276 326068 282328 326120
rect 309784 325592 309836 325644
rect 580172 325592 580224 325644
rect 266636 325388 266688 325440
rect 311900 325388 311952 325440
rect 268752 325320 268804 325372
rect 322940 325320 322992 325372
rect 276296 325252 276348 325304
rect 400220 325252 400272 325304
rect 292304 325184 292356 325236
rect 457444 325184 457496 325236
rect 115204 325116 115256 325168
rect 242256 325116 242308 325168
rect 286048 325116 286100 325168
rect 496820 325116 496872 325168
rect 107568 325048 107620 325100
rect 245936 325048 245988 325100
rect 252928 325048 252980 325100
rect 69664 324980 69716 325032
rect 242072 324980 242124 325032
rect 53748 324912 53800 324964
rect 240508 324912 240560 324964
rect 288164 325048 288216 325100
rect 510620 325048 510672 325100
rect 289544 324980 289596 325032
rect 524420 324980 524472 325032
rect 290832 324912 290884 324964
rect 542360 324912 542412 324964
rect 253020 324844 253072 324896
rect 268844 323892 268896 323944
rect 329840 323892 329892 323944
rect 276664 323824 276716 323876
rect 403624 323824 403676 323876
rect 293408 323756 293460 323808
rect 447784 323756 447836 323808
rect 291568 323688 291620 323740
rect 454684 323688 454736 323740
rect 286416 323620 286468 323672
rect 499580 323620 499632 323672
rect 234988 323595 235040 323604
rect 234988 323561 234997 323595
rect 234997 323561 235031 323595
rect 235031 323561 235040 323595
rect 234988 323552 235040 323561
rect 287244 323552 287296 323604
rect 514852 323552 514904 323604
rect 251364 323008 251416 323060
rect 251732 323008 251784 323060
rect 277032 322328 277084 322380
rect 407212 322328 407264 322380
rect 291936 322260 291988 322312
rect 483664 322260 483716 322312
rect 288900 322192 288952 322244
rect 528560 322192 528612 322244
rect 283932 321580 283984 321632
rect 284116 321580 284168 321632
rect 3516 320084 3568 320136
rect 234068 320084 234120 320136
rect 252928 319268 252980 319320
rect 253112 319268 253164 319320
rect 316684 313216 316736 313268
rect 580172 313216 580224 313268
rect 3516 306280 3568 306332
rect 209044 306280 209096 306332
rect 300216 299412 300268 299464
rect 580172 299412 580224 299464
rect 3056 293904 3108 293956
rect 222936 293904 222988 293956
rect 323676 289076 323728 289128
rect 512000 289076 512052 289128
rect 307116 273164 307168 273216
rect 580172 273164 580224 273216
rect 3516 267656 3568 267708
rect 232596 267656 232648 267708
rect 314016 259360 314068 259412
rect 580172 259360 580224 259412
rect 298836 245556 298888 245608
rect 580172 245556 580224 245608
rect 3516 241408 3568 241460
rect 220176 241408 220228 241460
rect 305644 233180 305696 233232
rect 579988 233180 580040 233232
rect 3332 215228 3384 215280
rect 231216 215228 231268 215280
rect 295984 206932 296036 206984
rect 579804 206932 579856 206984
rect 304264 193128 304316 193180
rect 580172 193128 580224 193180
rect 3516 188980 3568 189032
rect 215944 188980 215996 189032
rect 324964 177284 325016 177336
rect 518900 177284 518952 177336
rect 583116 165903 583168 165912
rect 583116 165869 583125 165903
rect 583125 165869 583159 165903
rect 583159 165869 583168 165903
rect 583116 165860 583168 165869
rect 2780 164092 2832 164144
rect 4804 164092 4856 164144
rect 583024 152711 583076 152720
rect 583024 152677 583033 152711
rect 583033 152677 583067 152711
rect 583067 152677 583076 152711
rect 583024 152668 583076 152677
rect 582840 126055 582892 126064
rect 582840 126021 582849 126055
rect 582849 126021 582883 126055
rect 582883 126021 582892 126055
rect 582840 126012 582892 126021
rect 582748 112863 582800 112872
rect 582748 112829 582757 112863
rect 582757 112829 582791 112863
rect 582791 112829 582800 112863
rect 582748 112820 582800 112829
rect 582656 99535 582708 99544
rect 582656 99501 582665 99535
rect 582665 99501 582699 99535
rect 582699 99501 582708 99535
rect 582656 99492 582708 99501
rect 582564 86207 582616 86216
rect 582564 86173 582573 86207
rect 582573 86173 582607 86207
rect 582607 86173 582616 86207
rect 582564 86164 582616 86173
rect 3148 85484 3200 85536
rect 214564 85484 214616 85536
rect 582472 73015 582524 73024
rect 582472 72981 582481 73015
rect 582481 72981 582515 73015
rect 582515 72981 582524 73015
rect 582472 72972 582524 72981
rect 3424 71680 3476 71732
rect 228456 71680 228508 71732
rect 582380 46359 582432 46368
rect 582380 46325 582389 46359
rect 582389 46325 582423 46359
rect 582423 46325 582432 46359
rect 582380 46316 582432 46325
rect 3424 45500 3476 45552
rect 213184 45500 213236 45552
rect 3148 33056 3200 33108
rect 226984 33056 227036 33108
rect 234712 33056 234764 33108
rect 580172 33056 580224 33108
rect 3424 20612 3476 20664
rect 294972 20612 295024 20664
rect 157248 17212 157300 17264
rect 250352 17212 250404 17264
rect 327724 17212 327776 17264
rect 550640 17212 550692 17264
rect 267188 15852 267240 15904
rect 316224 15852 316276 15904
rect 323584 15512 323636 15564
rect 328000 15512 328052 15564
rect 215208 14424 215260 14476
rect 222844 14424 222896 14476
rect 287612 13132 287664 13184
rect 517888 13132 517940 13184
rect 5264 13064 5316 13116
rect 173164 13064 173216 13116
rect 228732 13064 228784 13116
rect 233976 13064 234028 13116
rect 292028 13064 292080 13116
rect 556896 13064 556948 13116
rect 280712 12112 280764 12164
rect 442632 12112 442684 12164
rect 280620 12044 280672 12096
rect 445760 12044 445812 12096
rect 280528 11976 280580 12028
rect 448520 11976 448572 12028
rect 281908 11908 281960 11960
rect 453212 11908 453264 11960
rect 282000 11840 282052 11892
rect 456892 11840 456944 11892
rect 165528 11772 165580 11824
rect 224224 11772 224276 11824
rect 282184 11772 282236 11824
rect 459928 11772 459980 11824
rect 65432 11704 65484 11756
rect 240508 11704 240560 11756
rect 282092 11704 282144 11756
rect 463976 11704 464028 11756
rect 324412 11636 324464 11688
rect 325608 11636 325660 11688
rect 407212 11636 407264 11688
rect 408408 11636 408460 11688
rect 423772 11636 423824 11688
rect 424968 11636 425020 11688
rect 272708 10956 272760 11008
rect 367744 10956 367796 11008
rect 272616 10888 272668 10940
rect 371240 10888 371292 10940
rect 273996 10820 274048 10872
rect 374000 10820 374052 10872
rect 274180 10752 274232 10804
rect 378416 10752 378468 10804
rect 274088 10684 274140 10736
rect 382372 10684 382424 10736
rect 275468 10616 275520 10668
rect 385592 10616 385644 10668
rect 275376 10548 275428 10600
rect 389456 10548 389508 10600
rect 150348 10480 150400 10532
rect 250168 10480 250220 10532
rect 275652 10480 275704 10532
rect 392584 10480 392636 10532
rect 122748 10412 122800 10464
rect 247500 10412 247552 10464
rect 275284 10412 275336 10464
rect 396080 10412 396132 10464
rect 119804 10344 119856 10396
rect 247408 10344 247460 10396
rect 276572 10344 276624 10396
rect 400128 10344 400180 10396
rect 115848 10276 115900 10328
rect 246396 10276 246448 10328
rect 277124 10276 277176 10328
rect 403532 10276 403584 10328
rect 272524 10208 272576 10260
rect 364616 10208 364668 10260
rect 272800 10140 272852 10192
rect 360752 10140 360804 10192
rect 271144 10072 271196 10124
rect 357532 10072 357584 10124
rect 271420 10004 271472 10056
rect 353576 10004 353628 10056
rect 270592 9936 270644 9988
rect 350448 9936 350500 9988
rect 271328 9868 271380 9920
rect 346952 9868 347004 9920
rect 270040 9800 270092 9852
rect 342904 9800 342956 9852
rect 270132 9732 270184 9784
rect 339500 9732 339552 9784
rect 231032 9392 231084 9444
rect 257436 9392 257488 9444
rect 160100 9324 160152 9376
rect 251548 9324 251600 9376
rect 266084 9324 266136 9376
rect 297272 9324 297324 9376
rect 142436 9256 142488 9308
rect 249248 9256 249300 9308
rect 265992 9256 266044 9308
rect 300768 9256 300820 9308
rect 138848 9188 138900 9240
rect 248696 9188 248748 9240
rect 265900 9188 265952 9240
rect 304356 9188 304408 9240
rect 135260 9120 135312 9172
rect 248972 9120 249024 9172
rect 268476 9120 268528 9172
rect 326804 9120 326856 9172
rect 83280 9052 83332 9104
rect 243360 9052 243412 9104
rect 284484 9052 284536 9104
rect 489920 9052 489972 9104
rect 79692 8984 79744 9036
rect 243268 8984 243320 9036
rect 294788 8984 294840 9036
rect 573916 8984 573968 9036
rect 8760 8916 8812 8968
rect 235356 8916 235408 8968
rect 294696 8916 294748 8968
rect 577412 8916 577464 8968
rect 199108 8168 199160 8220
rect 255964 8168 256016 8220
rect 181444 8100 181496 8152
rect 252928 8100 252980 8152
rect 174268 8032 174320 8084
rect 253020 8032 253072 8084
rect 170772 7964 170824 8016
rect 251640 7964 251692 8016
rect 280988 7964 281040 8016
rect 441528 7964 441580 8016
rect 167184 7896 167236 7948
rect 252008 7896 252060 7948
rect 280896 7896 280948 7948
rect 445024 7896 445076 7948
rect 163688 7828 163740 7880
rect 251364 7828 251416 7880
rect 281080 7828 281132 7880
rect 448612 7828 448664 7880
rect 158904 7760 158956 7812
rect 251456 7760 251508 7812
rect 280804 7760 280856 7812
rect 452108 7760 452160 7812
rect 131764 7692 131816 7744
rect 248788 7692 248840 7744
rect 282276 7692 282328 7744
rect 455696 7692 455748 7744
rect 128176 7624 128228 7676
rect 247316 7624 247368 7676
rect 282460 7624 282512 7676
rect 459192 7624 459244 7676
rect 9956 7556 10008 7608
rect 177304 7556 177356 7608
rect 177856 7556 177908 7608
rect 253112 7556 253164 7608
rect 282368 7556 282420 7608
rect 462780 7556 462832 7608
rect 234620 6808 234672 6860
rect 580172 6808 580224 6860
rect 3332 6740 3384 6792
rect 294604 6740 294656 6792
rect 208584 6672 208636 6724
rect 255872 6672 255924 6724
rect 271604 6672 271656 6724
rect 356336 6672 356388 6724
rect 205088 6604 205140 6656
rect 255688 6604 255740 6656
rect 273076 6604 273128 6656
rect 359924 6604 359976 6656
rect 201500 6536 201552 6588
rect 255780 6536 255832 6588
rect 272984 6536 273036 6588
rect 363512 6536 363564 6588
rect 183744 6468 183796 6520
rect 252836 6468 252888 6520
rect 273168 6468 273220 6520
rect 367008 6468 367060 6520
rect 176660 6400 176712 6452
rect 253388 6400 253440 6452
rect 272892 6400 272944 6452
rect 370596 6400 370648 6452
rect 102232 6332 102284 6384
rect 180064 6332 180116 6384
rect 180248 6332 180300 6384
rect 253664 6332 253716 6384
rect 274272 6332 274324 6384
rect 374092 6332 374144 6384
rect 173164 6264 173216 6316
rect 252744 6264 252796 6316
rect 273720 6264 273772 6316
rect 377680 6264 377732 6316
rect 28816 6196 28868 6248
rect 130384 6196 130436 6248
rect 130568 6196 130620 6248
rect 247224 6196 247276 6248
rect 273904 6196 273956 6248
rect 381176 6196 381228 6248
rect 4068 6128 4120 6180
rect 235264 6128 235316 6180
rect 267004 6128 267056 6180
rect 273628 6128 273680 6180
rect 273812 6128 273864 6180
rect 384764 6128 384816 6180
rect 271512 6060 271564 6112
rect 352840 6060 352892 6112
rect 271052 5992 271104 6044
rect 349252 5992 349304 6044
rect 270960 5924 271012 5976
rect 345756 5924 345808 5976
rect 269856 5856 269908 5908
rect 342168 5856 342220 5908
rect 269948 5788 270000 5840
rect 338672 5788 338724 5840
rect 269672 5720 269724 5772
rect 335084 5720 335136 5772
rect 268660 5652 268712 5704
rect 331588 5652 331640 5704
rect 196808 5516 196860 5568
rect 202144 5516 202196 5568
rect 218060 5448 218112 5500
rect 232504 5448 232556 5500
rect 233056 5448 233108 5500
rect 253480 5448 253532 5500
rect 253848 5448 253900 5500
rect 267740 5448 267792 5500
rect 272432 5448 272484 5500
rect 284392 5448 284444 5500
rect 288992 5448 289044 5500
rect 289544 5448 289596 5500
rect 189724 5380 189776 5432
rect 233884 5380 233936 5432
rect 240508 5380 240560 5432
rect 258724 5380 258776 5432
rect 263140 5380 263192 5432
rect 276020 5380 276072 5432
rect 186136 5312 186188 5364
rect 204904 5312 204956 5364
rect 211068 5312 211120 5364
rect 255412 5312 255464 5364
rect 262496 5312 262548 5364
rect 278320 5312 278372 5364
rect 171968 5244 172020 5296
rect 206284 5244 206336 5296
rect 207388 5244 207440 5296
rect 255596 5244 255648 5296
rect 264428 5244 264480 5296
rect 279516 5244 279568 5296
rect 182548 5176 182600 5228
rect 196624 5176 196676 5228
rect 203892 5176 203944 5228
rect 256056 5176 256108 5228
rect 264520 5176 264572 5228
rect 281908 5176 281960 5228
rect 376116 5176 376168 5228
rect 402520 5176 402572 5228
rect 175464 5108 175516 5160
rect 198004 5108 198056 5160
rect 200304 5108 200356 5160
rect 255504 5108 255556 5160
rect 264336 5108 264388 5160
rect 283104 5108 283156 5160
rect 336004 5108 336056 5160
rect 391848 5108 391900 5160
rect 393964 5108 394016 5160
rect 409604 5108 409656 5160
rect 129372 5040 129424 5092
rect 247132 5040 247184 5092
rect 264612 5040 264664 5092
rect 285404 5040 285456 5092
rect 286324 5040 286376 5092
rect 309048 5040 309100 5092
rect 331864 5040 331916 5092
rect 495900 5040 495952 5092
rect 7656 4972 7708 5024
rect 2872 4904 2924 4956
rect 234620 4972 234672 5024
rect 254584 4972 254636 5024
rect 264704 4972 264756 5024
rect 286600 4972 286652 5024
rect 298744 4972 298796 5024
rect 235172 4904 235224 4956
rect 238116 4904 238168 4956
rect 258356 4904 258408 4956
rect 267280 4904 267332 4956
rect 319720 4904 319772 4956
rect 320824 4972 320876 5024
rect 494704 4972 494756 5024
rect 320916 4904 320968 4956
rect 322204 4904 322256 4956
rect 505376 4904 505428 4956
rect 1676 4836 1728 4888
rect 234896 4836 234948 4888
rect 239312 4836 239364 4888
rect 259736 4836 259788 4888
rect 264152 4836 264204 4888
rect 288992 4836 289044 4888
rect 289544 4836 289596 4888
rect 532516 4836 532568 4888
rect 572 4768 624 4820
rect 221556 4700 221608 4752
rect 231124 4700 231176 4752
rect 235080 4768 235132 4820
rect 237012 4768 237064 4820
rect 258632 4768 258684 4820
rect 265808 4768 265860 4820
rect 292580 4768 292632 4820
rect 294972 4768 295024 4820
rect 576308 4768 576360 4820
rect 234988 4700 235040 4752
rect 231676 4632 231728 4684
rect 249984 4700 250036 4752
rect 263048 4700 263100 4752
rect 274824 4700 274876 4752
rect 241704 4632 241756 4684
rect 258816 4632 258868 4684
rect 262956 4632 263008 4684
rect 271236 4632 271288 4684
rect 242900 4564 242952 4616
rect 259828 4564 259880 4616
rect 231768 4496 231820 4548
rect 247592 4496 247644 4548
rect 246396 4428 246448 4480
rect 259644 4428 259696 4480
rect 244096 4360 244148 4412
rect 251824 4360 251876 4412
rect 277124 4360 277176 4412
rect 277676 4360 277728 4412
rect 290188 4292 290240 4344
rect 295432 4292 295484 4344
rect 293684 4224 293736 4276
rect 295524 4224 295576 4276
rect 41880 4088 41932 4140
rect 83464 4088 83516 4140
rect 85672 4088 85724 4140
rect 193220 4156 193272 4208
rect 195244 4156 195296 4208
rect 225144 4156 225196 4208
rect 228364 4156 228416 4208
rect 234528 4156 234580 4208
rect 235816 4156 235868 4208
rect 280712 4156 280764 4208
rect 285680 4156 285732 4208
rect 289084 4156 289136 4208
rect 294880 4156 294932 4208
rect 497464 4156 497516 4208
rect 498200 4156 498252 4208
rect 499580 4156 499632 4208
rect 500592 4156 500644 4208
rect 522304 4156 522356 4208
rect 523040 4156 523092 4208
rect 60832 4020 60884 4072
rect 65432 4020 65484 4072
rect 78588 4020 78640 4072
rect 243176 4088 243228 4140
rect 257068 4088 257120 4140
rect 260104 4088 260156 4140
rect 281356 4088 281408 4140
rect 440332 4088 440384 4140
rect 453304 4088 453356 4140
rect 560852 4088 560904 4140
rect 52552 3952 52604 4004
rect 57244 3952 57296 4004
rect 82084 3952 82136 4004
rect 242992 4020 243044 4072
rect 251180 4020 251232 4072
rect 259920 4020 259972 4072
rect 281264 4020 281316 4072
rect 443644 4020 443696 4072
rect 571524 4020 571576 4072
rect 243452 3952 243504 4004
rect 281172 3952 281224 4004
rect 447416 3952 447468 4004
rect 44272 3884 44324 3936
rect 50344 3884 50396 3936
rect 64328 3884 64380 3936
rect 68376 3884 68428 3936
rect 75000 3884 75052 3936
rect 241980 3884 242032 3936
rect 248788 3884 248840 3936
rect 260196 3884 260248 3936
rect 281448 3884 281500 3936
rect 450084 3952 450136 4004
rect 450544 3952 450596 4004
rect 447784 3884 447836 3936
rect 568028 3952 568080 4004
rect 23020 3816 23072 3868
rect 43444 3816 43496 3868
rect 46664 3816 46716 3868
rect 239128 3816 239180 3868
rect 282828 3816 282880 3868
rect 564440 3884 564492 3936
rect 18236 3748 18288 3800
rect 39396 3748 39448 3800
rect 43076 3748 43128 3800
rect 39580 3680 39632 3732
rect 238024 3748 238076 3800
rect 255872 3748 255924 3800
rect 260932 3748 260984 3800
rect 282644 3748 282696 3800
rect 454500 3748 454552 3800
rect 454684 3748 454736 3800
rect 550272 3816 550324 3868
rect 457444 3748 457496 3800
rect 546684 3748 546736 3800
rect 32312 3612 32364 3664
rect 27712 3544 27764 3596
rect 28908 3544 28960 3596
rect 31300 3544 31352 3596
rect 32496 3544 32548 3596
rect 33600 3544 33652 3596
rect 34428 3544 34480 3596
rect 35992 3612 36044 3664
rect 239220 3680 239272 3732
rect 254676 3680 254728 3732
rect 261208 3680 261260 3732
rect 282736 3680 282788 3732
rect 461584 3680 461636 3732
rect 461676 3680 461728 3732
rect 239404 3612 239456 3664
rect 282552 3612 282604 3664
rect 465172 3612 465224 3664
rect 237840 3544 237892 3596
rect 252376 3544 252428 3596
rect 261024 3544 261076 3596
rect 263416 3544 263468 3596
rect 266544 3544 266596 3596
rect 283748 3544 283800 3596
rect 468668 3612 468720 3664
rect 539600 3612 539652 3664
rect 468484 3544 468536 3596
rect 469864 3544 469916 3596
rect 514760 3544 514812 3596
rect 515956 3544 516008 3596
rect 524420 3544 524472 3596
rect 525432 3544 525484 3596
rect 17040 3476 17092 3528
rect 17868 3476 17920 3528
rect 25320 3476 25372 3528
rect 13544 3408 13596 3460
rect 22744 3408 22796 3460
rect 24216 3408 24268 3460
rect 229836 3476 229888 3528
rect 230388 3476 230440 3528
rect 232228 3476 232280 3528
rect 233148 3476 233200 3528
rect 233424 3476 233476 3528
rect 234436 3476 234488 3528
rect 259460 3476 259512 3528
rect 261116 3476 261168 3528
rect 262128 3476 262180 3528
rect 262956 3476 263008 3528
rect 264244 3476 264296 3528
rect 265348 3476 265400 3528
rect 283932 3476 283984 3528
rect 472256 3476 472308 3528
rect 237656 3408 237708 3460
rect 245200 3408 245252 3460
rect 257344 3408 257396 3460
rect 262864 3408 262916 3460
rect 264152 3408 264204 3460
rect 284024 3408 284076 3460
rect 475752 3476 475804 3528
rect 510068 3476 510120 3528
rect 510712 3476 510764 3528
rect 512644 3476 512696 3528
rect 513564 3476 513616 3528
rect 519544 3476 519596 3528
rect 521844 3476 521896 3528
rect 530584 3476 530636 3528
rect 531320 3476 531372 3528
rect 534908 3476 534960 3528
rect 535460 3476 535512 3528
rect 541992 3476 542044 3528
rect 542452 3476 542504 3528
rect 545488 3476 545540 3528
rect 546500 3476 546552 3528
rect 551284 3476 551336 3528
rect 552664 3476 552716 3528
rect 559748 3476 559800 3528
rect 560300 3476 560352 3528
rect 472624 3408 472676 3460
rect 473452 3408 473504 3460
rect 483756 3408 483808 3460
rect 553768 3408 553820 3460
rect 566556 3408 566608 3460
rect 572720 3408 572772 3460
rect 26516 3340 26568 3392
rect 29644 3340 29696 3392
rect 30104 3340 30156 3392
rect 32404 3340 32456 3392
rect 34796 3340 34848 3392
rect 35808 3340 35860 3392
rect 38384 3340 38436 3392
rect 39304 3340 39356 3392
rect 40684 3340 40736 3392
rect 41328 3340 41380 3392
rect 50160 3340 50212 3392
rect 50988 3340 51040 3392
rect 51356 3340 51408 3392
rect 52368 3340 52420 3392
rect 56048 3340 56100 3392
rect 57336 3340 57388 3392
rect 58440 3340 58492 3392
rect 59268 3340 59320 3392
rect 59636 3340 59688 3392
rect 61384 3340 61436 3392
rect 65524 3340 65576 3392
rect 66168 3340 66220 3392
rect 66720 3340 66772 3392
rect 68284 3340 68336 3392
rect 69112 3340 69164 3392
rect 70216 3340 70268 3392
rect 70308 3340 70360 3392
rect 71044 3340 71096 3392
rect 72608 3340 72660 3392
rect 73068 3340 73120 3392
rect 76196 3340 76248 3392
rect 77208 3340 77260 3392
rect 77392 3340 77444 3392
rect 79324 3340 79376 3392
rect 80888 3340 80940 3392
rect 81348 3340 81400 3392
rect 90364 3340 90416 3392
rect 91008 3340 91060 3392
rect 91560 3340 91612 3392
rect 93124 3340 93176 3392
rect 93952 3340 94004 3392
rect 95056 3340 95108 3392
rect 97448 3340 97500 3392
rect 97908 3340 97960 3392
rect 98644 3340 98696 3392
rect 99288 3340 99340 3392
rect 101036 3340 101088 3392
rect 102048 3340 102100 3392
rect 67916 3272 67968 3324
rect 69664 3272 69716 3324
rect 87972 3272 88024 3324
rect 88984 3272 89036 3324
rect 11152 3204 11204 3256
rect 14464 3204 14516 3256
rect 57244 3204 57296 3256
rect 58624 3204 58676 3256
rect 89168 3204 89220 3256
rect 243084 3340 243136 3392
rect 279976 3340 280028 3392
rect 244556 3272 244608 3324
rect 279792 3272 279844 3324
rect 48964 3068 49016 3120
rect 53104 3068 53156 3120
rect 96252 3068 96304 3120
rect 244740 3204 244792 3256
rect 279884 3204 279936 3256
rect 425704 3272 425756 3324
rect 427268 3272 427320 3324
rect 432604 3340 432656 3392
rect 434444 3340 434496 3392
rect 436744 3340 436796 3392
rect 437940 3340 437992 3392
rect 448520 3340 448572 3392
rect 449808 3340 449860 3392
rect 458088 3340 458140 3392
rect 464344 3340 464396 3392
rect 536104 3340 536156 3392
rect 443828 3272 443880 3324
rect 244832 3136 244884 3188
rect 258264 3136 258316 3188
rect 261300 3136 261352 3188
rect 263508 3136 263560 3188
rect 270040 3136 270092 3188
rect 279608 3136 279660 3188
rect 103336 3068 103388 3120
rect 245108 3068 245160 3120
rect 278136 3068 278188 3120
rect 414664 3136 414716 3188
rect 416688 3136 416740 3188
rect 19432 3000 19484 3052
rect 25504 3000 25556 3052
rect 92756 3000 92808 3052
rect 105728 3000 105780 3052
rect 106188 3000 106240 3052
rect 106924 3000 106976 3052
rect 107568 3000 107620 3052
rect 108120 3000 108172 3052
rect 108948 3000 109000 3052
rect 109316 3000 109368 3052
rect 111064 3000 111116 3052
rect 111156 3000 111208 3052
rect 246212 3000 246264 3052
rect 263324 3000 263376 3052
rect 268844 3000 268896 3052
rect 277952 3000 278004 3052
rect 73804 2932 73856 2984
rect 75184 2932 75236 2984
rect 71504 2864 71556 2916
rect 115112 2932 115164 2984
rect 115204 2932 115256 2984
rect 115848 2932 115900 2984
rect 116400 2932 116452 2984
rect 117228 2932 117280 2984
rect 118792 2932 118844 2984
rect 119804 2932 119856 2984
rect 84476 2864 84528 2916
rect 87604 2864 87656 2916
rect 99840 2864 99892 2916
rect 114008 2864 114060 2916
rect 122104 2932 122156 2984
rect 122288 2932 122340 2984
rect 122748 2932 122800 2984
rect 123484 2932 123536 2984
rect 124128 2932 124180 2984
rect 124680 2932 124732 2984
rect 125416 2932 125468 2984
rect 125876 2932 125928 2984
rect 126888 2932 126940 2984
rect 126980 2932 127032 2984
rect 129004 2932 129056 2984
rect 246120 2932 246172 2984
rect 278504 2932 278556 2984
rect 121092 2864 121144 2916
rect 110512 2796 110564 2848
rect 111156 2796 111208 2848
rect 117596 2796 117648 2848
rect 247500 2864 247552 2916
rect 276756 2864 276808 2916
rect 132960 2796 133012 2848
rect 133788 2796 133840 2848
rect 134156 2796 134208 2848
rect 135168 2796 135220 2848
rect 136456 2796 136508 2848
rect 137284 2796 137336 2848
rect 140044 2796 140096 2848
rect 140688 2796 140740 2848
rect 141240 2796 141292 2848
rect 142068 2796 142120 2848
rect 143540 2796 143592 2848
rect 144828 2796 144880 2848
rect 147128 2796 147180 2848
rect 147588 2796 147640 2848
rect 148324 2796 148376 2848
rect 148968 2796 149020 2848
rect 149520 2796 149572 2848
rect 150348 2796 150400 2848
rect 150624 2796 150676 2848
rect 151728 2796 151780 2848
rect 151820 2796 151872 2848
rect 153108 2796 153160 2848
rect 154212 2796 154264 2848
rect 155224 2796 155276 2848
rect 155408 2796 155460 2848
rect 155868 2796 155920 2848
rect 156604 2796 156656 2848
rect 157248 2796 157300 2848
rect 157800 2796 157852 2848
rect 158628 2796 158680 2848
rect 164884 2796 164936 2848
rect 165528 2796 165580 2848
rect 166080 2796 166132 2848
rect 166908 2796 166960 2848
rect 168380 2796 168432 2848
rect 169668 2796 169720 2848
rect 188528 2796 188580 2848
rect 188988 2796 189040 2848
rect 190828 2796 190880 2848
rect 191748 2796 191800 2848
rect 192024 2796 192076 2848
rect 193128 2796 193180 2848
rect 197912 2796 197964 2848
rect 198648 2796 198700 2848
rect 206192 2796 206244 2848
rect 206928 2796 206980 2848
rect 209780 2796 209832 2848
rect 210976 2796 211028 2848
rect 213368 2796 213420 2848
rect 213828 2796 213880 2848
rect 214472 2796 214524 2848
rect 215208 2796 215260 2848
rect 215668 2796 215720 2848
rect 216588 2796 216640 2848
rect 216864 2796 216916 2848
rect 217968 2796 218020 2848
rect 219256 2796 219308 2848
rect 220084 2796 220136 2848
rect 222752 2796 222804 2848
rect 223488 2796 223540 2848
rect 223948 2796 224000 2848
rect 224868 2796 224920 2848
rect 226340 2796 226392 2848
rect 227444 2796 227496 2848
rect 237932 2796 237984 2848
rect 300124 2796 300176 2848
rect 301964 2796 302016 2848
rect 307024 2796 307076 2848
rect 307944 2796 307996 2848
rect 313924 2796 313976 2848
rect 315028 2796 315080 2848
rect 316040 2796 316092 2848
rect 317328 2796 317380 2848
rect 331956 2796 332008 2848
rect 332692 2796 332744 2848
rect 333980 2796 334032 2848
rect 337476 2796 337528 2848
rect 338120 2796 338172 2848
rect 342996 2796 343048 2848
rect 344560 2796 344612 2848
rect 348056 2796 348108 2848
rect 349160 2796 349212 2848
rect 353944 2796 353996 2848
rect 355232 2796 355284 2848
rect 357440 2796 357492 2848
rect 358728 2796 358780 2848
rect 360844 2796 360896 2848
rect 362316 2796 362368 2848
rect 365812 2796 365864 2848
rect 367100 2796 367152 2848
rect 369400 2796 369452 2848
rect 369860 2796 369912 2848
rect 371884 2796 371936 2848
rect 372896 2796 372948 2848
rect 374000 2796 374052 2848
rect 375288 2796 375340 2848
rect 378784 2796 378836 2848
rect 379980 2796 380032 2848
rect 382280 2796 382332 2848
rect 383568 2796 383620 2848
rect 385684 2796 385736 2848
rect 387156 2796 387208 2848
rect 389824 2796 389876 2848
rect 390652 2796 390704 2848
rect 392676 2796 392728 2848
rect 394240 2796 394292 2848
rect 396724 2864 396776 2916
rect 397736 2864 397788 2916
rect 403624 2864 403676 2916
rect 404820 2864 404872 2916
rect 415492 3000 415544 3052
rect 418804 3068 418856 3120
rect 420184 3068 420236 3120
rect 433248 3204 433300 3256
rect 436744 3204 436796 3256
rect 490564 3204 490616 3256
rect 492312 3204 492364 3256
rect 578608 3204 578660 3256
rect 560944 3136 560996 3188
rect 563244 3136 563296 3188
rect 429660 3068 429712 3120
rect 426164 3000 426216 3052
rect 527824 3000 527876 3052
rect 528652 3000 528704 3052
rect 422576 2932 422628 2984
rect 411904 2796 411956 2848
rect 418988 2796 419040 2848
rect 450084 2796 450136 2848
rect 450912 2796 450964 2848
rect 333888 2728 333940 2780
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 89364 703582 89668 703610
rect 8128 700534 8156 703520
rect 8116 700528 8168 700534
rect 8116 700470 8168 700476
rect 24320 699718 24348 703520
rect 40512 700398 40540 703520
rect 72988 700806 73016 703520
rect 89180 703474 89208 703520
rect 89364 703474 89392 703582
rect 89180 703446 89392 703474
rect 72976 700800 73028 700806
rect 72976 700742 73028 700748
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 41328 700392 41380 700398
rect 41328 700334 41380 700340
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3146 658200 3202 658209
rect 3146 658135 3202 658144
rect 3160 656946 3188 658135
rect 3148 656940 3200 656946
rect 3148 656882 3200 656888
rect 3330 606112 3386 606121
rect 3330 606047 3386 606056
rect 3344 605878 3372 606047
rect 3332 605872 3384 605878
rect 3332 605814 3384 605820
rect 3146 553888 3202 553897
rect 3146 553823 3202 553832
rect 3160 553450 3188 553823
rect 3148 553444 3200 553450
rect 3148 553386 3200 553392
rect 3238 501800 3294 501809
rect 3238 501735 3294 501744
rect 3252 501022 3280 501735
rect 3240 501016 3292 501022
rect 3240 500958 3292 500964
rect 3330 475688 3386 475697
rect 3330 475623 3386 475632
rect 3238 462632 3294 462641
rect 3238 462567 3294 462576
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 3146 423600 3202 423609
rect 3146 423535 3202 423544
rect 3054 410544 3110 410553
rect 3054 410479 3110 410488
rect 2964 397520 3016 397526
rect 2962 397488 2964 397497
rect 3016 397488 3018 397497
rect 2962 397423 3018 397432
rect 3068 380186 3096 410479
rect 3160 380254 3188 423535
rect 3252 380322 3280 462567
rect 3344 380390 3372 475623
rect 3332 380384 3384 380390
rect 3332 380326 3384 380332
rect 3240 380316 3292 380322
rect 3240 380258 3292 380264
rect 3148 380248 3200 380254
rect 3436 380225 3464 684247
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 380798 3556 671191
rect 3606 632088 3662 632097
rect 3606 632023 3662 632032
rect 3620 380866 3648 632023
rect 3698 619168 3754 619177
rect 3698 619103 3754 619112
rect 3608 380860 3660 380866
rect 3608 380802 3660 380808
rect 3516 380792 3568 380798
rect 3516 380734 3568 380740
rect 3712 380730 3740 619103
rect 3790 580000 3846 580009
rect 3790 579935 3846 579944
rect 3700 380724 3752 380730
rect 3700 380666 3752 380672
rect 3804 380594 3832 579935
rect 3882 566944 3938 566953
rect 3882 566879 3938 566888
rect 3896 380662 3924 566879
rect 3974 527912 4030 527921
rect 3974 527847 4030 527856
rect 3884 380656 3936 380662
rect 3884 380598 3936 380604
rect 3792 380588 3844 380594
rect 3792 380530 3844 380536
rect 3988 380526 4016 527847
rect 4066 514856 4122 514865
rect 4066 514791 4122 514800
rect 3976 380520 4028 380526
rect 3976 380462 4028 380468
rect 4080 380458 4108 514791
rect 4068 380452 4120 380458
rect 4068 380394 4120 380400
rect 24780 380361 24808 699654
rect 24766 380352 24822 380361
rect 24766 380287 24822 380296
rect 3148 380190 3200 380196
rect 3422 380216 3478 380225
rect 3056 380180 3108 380186
rect 3422 380151 3478 380160
rect 3056 380122 3108 380128
rect 41340 380118 41368 700334
rect 41328 380112 41380 380118
rect 41328 380054 41380 380060
rect 89640 379982 89668 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 154316 703582 154528 703610
rect 105464 699718 105492 703520
rect 137848 700262 137876 703520
rect 154132 703474 154160 703520
rect 154316 703474 154344 703582
rect 154132 703446 154344 703474
rect 137836 700256 137888 700262
rect 137836 700198 137888 700204
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 106200 380050 106228 699654
rect 106188 380044 106240 380050
rect 106188 379986 106240 379992
rect 89628 379976 89680 379982
rect 89628 379918 89680 379924
rect 154500 379914 154528 703582
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 170324 699718 170352 703520
rect 202800 699990 202828 703520
rect 218992 702434 219020 703520
rect 218992 702406 219388 702434
rect 202788 699984 202840 699990
rect 202788 699926 202840 699932
rect 170312 699712 170364 699718
rect 170312 699654 170364 699660
rect 171048 699712 171100 699718
rect 171048 699654 171100 699660
rect 154488 379908 154540 379914
rect 154488 379850 154540 379856
rect 171060 379846 171088 699654
rect 171048 379840 171100 379846
rect 171048 379782 171100 379788
rect 219360 379778 219388 702406
rect 235184 699718 235212 703520
rect 263324 701004 263376 701010
rect 263324 700946 263376 700952
rect 262036 700868 262088 700874
rect 262036 700810 262088 700816
rect 261944 700664 261996 700670
rect 261944 700606 261996 700612
rect 260656 700596 260708 700602
rect 260656 700538 260708 700544
rect 259368 700460 259420 700466
rect 259368 700402 259420 700408
rect 259276 700324 259328 700330
rect 259276 700266 259328 700272
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 235908 699712 235960 699718
rect 235908 699654 235960 699660
rect 219348 379772 219400 379778
rect 219348 379714 219400 379720
rect 235920 379642 235948 699654
rect 257988 696992 258040 696998
rect 257988 696934 258040 696940
rect 257896 670744 257948 670750
rect 257896 670686 257948 670692
rect 256608 643136 256660 643142
rect 256608 643078 256660 643084
rect 256516 616888 256568 616894
rect 256516 616830 256568 616836
rect 255228 590708 255280 590714
rect 255228 590650 255280 590656
rect 255136 576904 255188 576910
rect 255136 576846 255188 576852
rect 255044 563100 255096 563106
rect 255044 563042 255096 563048
rect 253848 536852 253900 536858
rect 253848 536794 253900 536800
rect 253756 524476 253808 524482
rect 253756 524418 253808 524424
rect 252468 510672 252520 510678
rect 252468 510614 252520 510620
rect 252376 484424 252428 484430
rect 252376 484366 252428 484372
rect 252284 470620 252336 470626
rect 252284 470562 252336 470568
rect 251088 456816 251140 456822
rect 251088 456758 251140 456764
rect 250996 430636 251048 430642
rect 250996 430578 251048 430584
rect 250904 418192 250956 418198
rect 250904 418134 250956 418140
rect 249708 404388 249760 404394
rect 249708 404330 249760 404336
rect 235908 379636 235960 379642
rect 235908 379578 235960 379584
rect 234068 379432 234120 379438
rect 234068 379374 234120 379380
rect 232596 379296 232648 379302
rect 232596 379238 232648 379244
rect 231216 379228 231268 379234
rect 231216 379170 231268 379176
rect 222936 379092 222988 379098
rect 222936 379034 222988 379040
rect 215944 378684 215996 378690
rect 215944 378626 215996 378632
rect 213184 378616 213236 378622
rect 213184 378558 213236 378564
rect 3608 378548 3660 378554
rect 3608 378490 3660 378496
rect 3516 377528 3568 377534
rect 3516 377470 3568 377476
rect 3424 377460 3476 377466
rect 3424 377402 3476 377408
rect 3148 346384 3200 346390
rect 3148 346326 3200 346332
rect 3160 345409 3188 346326
rect 3146 345400 3202 345409
rect 3146 345335 3202 345344
rect 3056 293956 3108 293962
rect 3056 293898 3108 293904
rect 3068 293185 3096 293898
rect 3054 293176 3110 293185
rect 3054 293111 3110 293120
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 2780 164144 2832 164150
rect 2780 164086 2832 164092
rect 2792 162897 2820 164086
rect 2778 162888 2834 162897
rect 2778 162823 2834 162832
rect 3436 110673 3464 377402
rect 3528 358465 3556 377470
rect 3620 371385 3648 378490
rect 209044 377120 209096 377126
rect 209044 377062 209096 377068
rect 4804 377052 4856 377058
rect 4804 376994 4856 377000
rect 3606 371376 3662 371385
rect 3606 371311 3662 371320
rect 3514 358456 3570 358465
rect 3514 358391 3570 358400
rect 3516 320136 3568 320142
rect 3516 320078 3568 320084
rect 3528 319297 3556 320078
rect 3514 319288 3570 319297
rect 3514 319223 3570 319232
rect 3516 306332 3568 306338
rect 3516 306274 3568 306280
rect 3528 306241 3556 306274
rect 3514 306232 3570 306241
rect 3514 306167 3570 306176
rect 3516 267708 3568 267714
rect 3516 267650 3568 267656
rect 3528 267209 3556 267650
rect 3514 267200 3570 267209
rect 3514 267135 3570 267144
rect 3514 255232 3570 255241
rect 3514 255167 3570 255176
rect 3528 254153 3556 255167
rect 3514 254144 3570 254153
rect 3514 254079 3570 254088
rect 3516 241460 3568 241466
rect 3516 241402 3568 241408
rect 3528 241097 3556 241402
rect 3514 241088 3570 241097
rect 3514 241023 3570 241032
rect 3514 202872 3570 202881
rect 3514 202807 3570 202816
rect 3528 201929 3556 202807
rect 3514 201920 3570 201929
rect 3514 201855 3570 201864
rect 3516 189032 3568 189038
rect 3516 188974 3568 188980
rect 3528 188873 3556 188974
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 4816 164150 4844 376994
rect 125508 337680 125560 337686
rect 125508 337622 125560 337628
rect 122104 337612 122156 337618
rect 122104 337554 122156 337560
rect 97908 337544 97960 337550
rect 97908 337486 97960 337492
rect 91008 337476 91060 337482
rect 91008 337418 91060 337424
rect 86868 337408 86920 337414
rect 86868 337350 86920 337356
rect 81348 337340 81400 337346
rect 81348 337282 81400 337288
rect 70308 337272 70360 337278
rect 70308 337214 70360 337220
rect 66168 337204 66220 337210
rect 66168 337146 66220 337152
rect 50344 337136 50396 337142
rect 50344 337078 50396 337084
rect 48228 337068 48280 337074
rect 48228 337010 48280 337016
rect 41328 337000 41380 337006
rect 41328 336942 41380 336948
rect 34428 336932 34480 336938
rect 34428 336874 34480 336880
rect 29644 336864 29696 336870
rect 29644 336806 29696 336812
rect 12348 336796 12400 336802
rect 12348 336738 12400 336744
rect 4804 164144 4856 164150
rect 4804 164086 4856 164092
rect 3514 138000 3570 138009
rect 3514 137935 3570 137944
rect 3528 136785 3556 137935
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3330 59256 3386 59265
rect 3330 59191 3386 59200
rect 3344 58585 3372 59191
rect 3330 58576 3386 58585
rect 3330 58511 3386 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3148 33108 3200 33114
rect 3148 33050 3200 33056
rect 3160 32473 3188 33050
rect 3146 32464 3202 32473
rect 3146 32399 3202 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 5264 13116 5316 13122
rect 5264 13058 5316 13064
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 3344 6497 3372 6734
rect 3330 6488 3386 6497
rect 3330 6423 3386 6432
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 2872 4956 2924 4962
rect 2872 4898 2924 4904
rect 1676 4888 1728 4894
rect 1676 4830 1728 4836
rect 572 4820 624 4826
rect 572 4762 624 4768
rect 584 480 612 4762
rect 1688 480 1716 4830
rect 2884 480 2912 4898
rect 4080 480 4108 6122
rect 5276 480 5304 13058
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 6458 3360 6514 3369
rect 6458 3295 6514 3304
rect 6472 480 6500 3295
rect 7668 480 7696 4966
rect 8772 480 8800 8910
rect 9956 7608 10008 7614
rect 9956 7550 10008 7556
rect 9968 480 9996 7550
rect 11152 3256 11204 3262
rect 11152 3198 11204 3204
rect 11164 480 11192 3198
rect 12360 480 12388 336738
rect 25502 336152 25558 336161
rect 25502 336087 25558 336096
rect 14462 336016 14518 336025
rect 14462 335951 14518 335960
rect 13544 3460 13596 3466
rect 13544 3402 13596 3408
rect 13556 480 13584 3402
rect 14476 3262 14504 335951
rect 17868 334620 17920 334626
rect 17868 334562 17920 334568
rect 15934 3632 15990 3641
rect 15934 3567 15990 3576
rect 14738 3496 14794 3505
rect 14738 3431 14794 3440
rect 14464 3256 14516 3262
rect 14464 3198 14516 3204
rect 14752 480 14780 3431
rect 15948 480 15976 3567
rect 17880 3534 17908 334562
rect 22008 333260 22060 333266
rect 22008 333202 22060 333208
rect 22020 6914 22048 333202
rect 22744 330540 22796 330546
rect 22744 330482 22796 330488
rect 21836 6886 22048 6914
rect 18236 3800 18288 3806
rect 18236 3742 18288 3748
rect 20626 3768 20682 3777
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 17052 480 17080 3470
rect 18248 480 18276 3742
rect 20626 3703 20682 3712
rect 19432 3052 19484 3058
rect 19432 2994 19484 3000
rect 19444 480 19472 2994
rect 20640 480 20668 3703
rect 21836 480 21864 6886
rect 22756 3466 22784 330482
rect 23020 3868 23072 3874
rect 23020 3810 23072 3816
rect 22744 3460 22796 3466
rect 22744 3402 22796 3408
rect 23032 480 23060 3810
rect 25320 3528 25372 3534
rect 25320 3470 25372 3476
rect 24216 3460 24268 3466
rect 24216 3402 24268 3408
rect 24228 480 24256 3402
rect 25332 480 25360 3470
rect 25516 3058 25544 336087
rect 28908 327752 28960 327758
rect 28908 327694 28960 327700
rect 28816 6248 28868 6254
rect 28816 6190 28868 6196
rect 27712 3596 27764 3602
rect 27712 3538 27764 3544
rect 26516 3392 26568 3398
rect 26516 3334 26568 3340
rect 25504 3052 25556 3058
rect 25504 2994 25556 3000
rect 26528 480 26556 3334
rect 27724 480 27752 3538
rect 28828 3210 28856 6190
rect 28920 3602 28948 327694
rect 28908 3596 28960 3602
rect 28908 3538 28960 3544
rect 29656 3398 29684 336806
rect 32404 331900 32456 331906
rect 32404 331842 32456 331848
rect 32312 3664 32364 3670
rect 32312 3606 32364 3612
rect 31300 3596 31352 3602
rect 31300 3538 31352 3544
rect 29644 3392 29696 3398
rect 29644 3334 29696 3340
rect 30104 3392 30156 3398
rect 30104 3334 30156 3340
rect 28828 3182 28948 3210
rect 28920 480 28948 3182
rect 30116 480 30144 3334
rect 31312 480 31340 3538
rect 32324 1850 32352 3606
rect 32416 3398 32444 331842
rect 32496 329112 32548 329118
rect 32496 329054 32548 329060
rect 32508 3602 32536 329054
rect 34440 3602 34468 336874
rect 39304 330676 39356 330682
rect 39304 330618 39356 330624
rect 37188 330608 37240 330614
rect 37188 330550 37240 330556
rect 35808 326392 35860 326398
rect 35808 326334 35860 326340
rect 32496 3596 32548 3602
rect 32496 3538 32548 3544
rect 33600 3596 33652 3602
rect 33600 3538 33652 3544
rect 34428 3596 34480 3602
rect 34428 3538 34480 3544
rect 32404 3392 32456 3398
rect 32404 3334 32456 3340
rect 32324 1822 32444 1850
rect 32416 480 32444 1822
rect 33612 480 33640 3538
rect 35820 3398 35848 326334
rect 35992 3664 36044 3670
rect 35992 3606 36044 3612
rect 34796 3392 34848 3398
rect 34796 3334 34848 3340
rect 35808 3392 35860 3398
rect 35808 3334 35860 3340
rect 34808 480 34836 3334
rect 36004 480 36032 3606
rect 37200 480 37228 330550
rect 39316 3398 39344 330618
rect 39396 329180 39448 329186
rect 39396 329122 39448 329128
rect 39408 3806 39436 329122
rect 39396 3800 39448 3806
rect 39396 3742 39448 3748
rect 39580 3732 39632 3738
rect 39580 3674 39632 3680
rect 38384 3392 38436 3398
rect 38384 3334 38436 3340
rect 39304 3392 39356 3398
rect 39304 3334 39356 3340
rect 38396 480 38424 3334
rect 39592 480 39620 3674
rect 41340 3398 41368 336942
rect 43444 327888 43496 327894
rect 43444 327830 43496 327836
rect 41880 4140 41932 4146
rect 41880 4082 41932 4088
rect 40684 3392 40736 3398
rect 40684 3334 40736 3340
rect 41328 3392 41380 3398
rect 41328 3334 41380 3340
rect 40696 480 40724 3334
rect 41892 480 41920 4082
rect 43456 3874 43484 327830
rect 45468 327820 45520 327826
rect 45468 327762 45520 327768
rect 44272 3936 44324 3942
rect 44272 3878 44324 3884
rect 43444 3868 43496 3874
rect 43444 3810 43496 3816
rect 43076 3800 43128 3806
rect 43076 3742 43128 3748
rect 43088 480 43116 3742
rect 44284 480 44312 3878
rect 45480 480 45508 327762
rect 48240 6914 48268 337010
rect 47872 6886 48268 6914
rect 46664 3868 46716 3874
rect 46664 3810 46716 3816
rect 46676 480 46704 3810
rect 47872 480 47900 6886
rect 50356 3942 50384 337078
rect 52368 334688 52420 334694
rect 52368 334630 52420 334636
rect 50988 326460 51040 326466
rect 50988 326402 51040 326408
rect 50344 3936 50396 3942
rect 50344 3878 50396 3884
rect 51000 3398 51028 326402
rect 52380 3398 52408 334630
rect 59268 333396 59320 333402
rect 59268 333338 59320 333344
rect 55128 333328 55180 333334
rect 55128 333270 55180 333276
rect 53104 331968 53156 331974
rect 53104 331910 53156 331916
rect 52552 4004 52604 4010
rect 52552 3946 52604 3952
rect 50160 3392 50212 3398
rect 50160 3334 50212 3340
rect 50988 3392 51040 3398
rect 50988 3334 51040 3340
rect 51356 3392 51408 3398
rect 51356 3334 51408 3340
rect 52368 3392 52420 3398
rect 52368 3334 52420 3340
rect 48964 3120 49016 3126
rect 48964 3062 49016 3068
rect 48976 480 49004 3062
rect 50172 480 50200 3334
rect 51368 480 51396 3334
rect 52564 480 52592 3946
rect 53116 3126 53144 331910
rect 53748 324964 53800 324970
rect 53748 324906 53800 324912
rect 53104 3120 53156 3126
rect 53104 3062 53156 3068
rect 53760 480 53788 324906
rect 55140 6914 55168 333270
rect 57244 330744 57296 330750
rect 57244 330686 57296 330692
rect 54956 6886 55168 6914
rect 54956 480 54984 6886
rect 57256 4010 57284 330686
rect 57336 329248 57388 329254
rect 57336 329190 57388 329196
rect 57244 4004 57296 4010
rect 57244 3946 57296 3952
rect 57348 3398 57376 329190
rect 58624 326528 58676 326534
rect 58624 326470 58676 326476
rect 56048 3392 56100 3398
rect 56048 3334 56100 3340
rect 57336 3392 57388 3398
rect 57336 3334 57388 3340
rect 58440 3392 58492 3398
rect 58440 3334 58492 3340
rect 56060 480 56088 3334
rect 57244 3256 57296 3262
rect 57244 3198 57296 3204
rect 57256 480 57284 3198
rect 58452 480 58480 3334
rect 58636 3262 58664 326470
rect 59280 3398 59308 333338
rect 62028 332036 62080 332042
rect 62028 331978 62080 331984
rect 61384 329316 61436 329322
rect 61384 329258 61436 329264
rect 60832 4072 60884 4078
rect 60832 4014 60884 4020
rect 59268 3392 59320 3398
rect 59268 3334 59320 3340
rect 59636 3392 59688 3398
rect 59636 3334 59688 3340
rect 58624 3256 58676 3262
rect 58624 3198 58676 3204
rect 59648 480 59676 3334
rect 60844 480 60872 4014
rect 61396 3398 61424 329258
rect 61384 3392 61436 3398
rect 61384 3334 61436 3340
rect 62040 480 62068 331978
rect 63408 329384 63460 329390
rect 63408 329326 63460 329332
rect 63420 6914 63448 329326
rect 65432 11756 65484 11762
rect 65432 11698 65484 11704
rect 63236 6886 63448 6914
rect 63236 480 63264 6886
rect 65444 4078 65472 11698
rect 65432 4072 65484 4078
rect 65432 4014 65484 4020
rect 64328 3936 64380 3942
rect 64328 3878 64380 3884
rect 64340 480 64368 3878
rect 66180 3398 66208 337146
rect 68284 330812 68336 330818
rect 68284 330754 68336 330760
rect 68296 3398 68324 330754
rect 68376 326596 68428 326602
rect 68376 326538 68428 326544
rect 68388 3942 68416 326538
rect 69664 325032 69716 325038
rect 69664 324974 69716 324980
rect 68376 3936 68428 3942
rect 68376 3878 68428 3884
rect 65524 3392 65576 3398
rect 65524 3334 65576 3340
rect 66168 3392 66220 3398
rect 66168 3334 66220 3340
rect 66720 3392 66772 3398
rect 66720 3334 66772 3340
rect 68284 3392 68336 3398
rect 68284 3334 68336 3340
rect 69112 3392 69164 3398
rect 69112 3334 69164 3340
rect 65536 480 65564 3334
rect 66732 480 66760 3334
rect 67916 3324 67968 3330
rect 67916 3266 67968 3272
rect 67928 480 67956 3266
rect 69124 480 69152 3334
rect 69676 3330 69704 324974
rect 70320 6914 70348 337214
rect 73068 333464 73120 333470
rect 73068 333406 73120 333412
rect 71044 329452 71096 329458
rect 71044 329394 71096 329400
rect 70228 6886 70348 6914
rect 70228 3398 70256 6886
rect 71056 3398 71084 329394
rect 73080 3398 73108 333406
rect 77208 332104 77260 332110
rect 77208 332046 77260 332052
rect 75184 329520 75236 329526
rect 75184 329462 75236 329468
rect 75000 3936 75052 3942
rect 75000 3878 75052 3884
rect 70216 3392 70268 3398
rect 70216 3334 70268 3340
rect 70308 3392 70360 3398
rect 70308 3334 70360 3340
rect 71044 3392 71096 3398
rect 71044 3334 71096 3340
rect 72608 3392 72660 3398
rect 72608 3334 72660 3340
rect 73068 3392 73120 3398
rect 73068 3334 73120 3340
rect 69664 3324 69716 3330
rect 69664 3266 69716 3272
rect 70320 480 70348 3334
rect 71504 2916 71556 2922
rect 71504 2858 71556 2864
rect 71516 480 71544 2858
rect 72620 480 72648 3334
rect 73804 2984 73856 2990
rect 73804 2926 73856 2932
rect 73816 480 73844 2926
rect 75012 480 75040 3878
rect 75196 2990 75224 329462
rect 77220 3398 77248 332046
rect 79324 330880 79376 330886
rect 79324 330822 79376 330828
rect 78588 4072 78640 4078
rect 78588 4014 78640 4020
rect 76196 3392 76248 3398
rect 76196 3334 76248 3340
rect 77208 3392 77260 3398
rect 77208 3334 77260 3340
rect 77392 3392 77444 3398
rect 77392 3334 77444 3340
rect 75184 2984 75236 2990
rect 75184 2926 75236 2932
rect 76208 480 76236 3334
rect 77404 480 77432 3334
rect 78600 480 78628 4014
rect 79336 3398 79364 330822
rect 79692 9036 79744 9042
rect 79692 8978 79744 8984
rect 79324 3392 79376 3398
rect 79324 3334 79376 3340
rect 79704 480 79732 8978
rect 81360 3398 81388 337282
rect 83464 333532 83516 333538
rect 83464 333474 83516 333480
rect 83280 9104 83332 9110
rect 83280 9046 83332 9052
rect 82084 4004 82136 4010
rect 82084 3946 82136 3952
rect 80888 3392 80940 3398
rect 80888 3334 80940 3340
rect 81348 3392 81400 3398
rect 81348 3334 81400 3340
rect 80900 480 80928 3334
rect 82096 480 82124 3946
rect 83292 480 83320 9046
rect 83476 4146 83504 333474
rect 83464 4140 83516 4146
rect 83464 4082 83516 4088
rect 85672 4140 85724 4146
rect 85672 4082 85724 4088
rect 84476 2916 84528 2922
rect 84476 2858 84528 2864
rect 84488 480 84516 2858
rect 85684 480 85712 4082
rect 86880 480 86908 337350
rect 87604 334756 87656 334762
rect 87604 334698 87656 334704
rect 87616 2922 87644 334698
rect 88984 333600 89036 333606
rect 88984 333542 89036 333548
rect 88996 3330 89024 333542
rect 91020 3398 91048 337418
rect 95148 332172 95200 332178
rect 95148 332114 95200 332120
rect 93124 329588 93176 329594
rect 93124 329530 93176 329536
rect 93136 3398 93164 329530
rect 95056 327956 95108 327962
rect 95056 327898 95108 327904
rect 95068 16574 95096 327898
rect 94976 16546 95096 16574
rect 90364 3392 90416 3398
rect 90364 3334 90416 3340
rect 91008 3392 91060 3398
rect 91008 3334 91060 3340
rect 91560 3392 91612 3398
rect 91560 3334 91612 3340
rect 93124 3392 93176 3398
rect 93124 3334 93176 3340
rect 93952 3392 94004 3398
rect 93952 3334 94004 3340
rect 87972 3324 88024 3330
rect 87972 3266 88024 3272
rect 88984 3324 89036 3330
rect 88984 3266 89036 3272
rect 87604 2916 87656 2922
rect 87604 2858 87656 2864
rect 87984 480 88012 3266
rect 89168 3256 89220 3262
rect 89168 3198 89220 3204
rect 89180 480 89208 3198
rect 90376 480 90404 3334
rect 91572 480 91600 3334
rect 92756 3052 92808 3058
rect 92756 2994 92808 3000
rect 92768 480 92796 2994
rect 93964 480 93992 3334
rect 94976 3210 95004 16546
rect 95160 6914 95188 332114
rect 95068 6886 95188 6914
rect 95068 3398 95096 6886
rect 97920 3398 97948 337486
rect 104808 332240 104860 332246
rect 104808 332182 104860 332188
rect 102048 330948 102100 330954
rect 102048 330890 102100 330896
rect 99288 329656 99340 329662
rect 99288 329598 99340 329604
rect 99300 3398 99328 329598
rect 102060 3398 102088 330890
rect 104820 6914 104848 332182
rect 111708 331084 111760 331090
rect 111708 331026 111760 331032
rect 108948 331016 109000 331022
rect 108948 330958 109000 330964
rect 106188 328024 106240 328030
rect 106188 327966 106240 327972
rect 104544 6886 104848 6914
rect 102232 6384 102284 6390
rect 102232 6326 102284 6332
rect 95056 3392 95108 3398
rect 95056 3334 95108 3340
rect 97448 3392 97500 3398
rect 97448 3334 97500 3340
rect 97908 3392 97960 3398
rect 97908 3334 97960 3340
rect 98644 3392 98696 3398
rect 98644 3334 98696 3340
rect 99288 3392 99340 3398
rect 99288 3334 99340 3340
rect 101036 3392 101088 3398
rect 101036 3334 101088 3340
rect 102048 3392 102100 3398
rect 102048 3334 102100 3340
rect 94976 3182 95188 3210
rect 95160 480 95188 3182
rect 96252 3120 96304 3126
rect 96252 3062 96304 3068
rect 96264 480 96292 3062
rect 97460 480 97488 3334
rect 98656 480 98684 3334
rect 99840 2916 99892 2922
rect 99840 2858 99892 2864
rect 99852 480 99880 2858
rect 101048 480 101076 3334
rect 102244 480 102272 6326
rect 103336 3120 103388 3126
rect 103336 3062 103388 3068
rect 103348 480 103376 3062
rect 104544 480 104572 6886
rect 106200 3058 106228 327966
rect 107568 325100 107620 325106
rect 107568 325042 107620 325048
rect 107580 3058 107608 325042
rect 108960 3058 108988 330958
rect 111064 328092 111116 328098
rect 111064 328034 111116 328040
rect 111076 3058 111104 328034
rect 111720 6914 111748 331026
rect 119988 328228 120040 328234
rect 119988 328170 120040 328176
rect 113088 328160 113140 328166
rect 113088 328102 113140 328108
rect 113100 6914 113128 328102
rect 117228 326664 117280 326670
rect 117228 326606 117280 326612
rect 115204 325168 115256 325174
rect 115204 325110 115256 325116
rect 115216 6914 115244 325110
rect 115848 10328 115900 10334
rect 115848 10270 115900 10276
rect 111628 6886 111748 6914
rect 112824 6886 113128 6914
rect 115124 6886 115244 6914
rect 105728 3052 105780 3058
rect 105728 2994 105780 3000
rect 106188 3052 106240 3058
rect 106188 2994 106240 3000
rect 106924 3052 106976 3058
rect 106924 2994 106976 3000
rect 107568 3052 107620 3058
rect 107568 2994 107620 3000
rect 108120 3052 108172 3058
rect 108120 2994 108172 3000
rect 108948 3052 109000 3058
rect 108948 2994 109000 3000
rect 109316 3052 109368 3058
rect 109316 2994 109368 3000
rect 111064 3052 111116 3058
rect 111064 2994 111116 3000
rect 111156 3052 111208 3058
rect 111156 2994 111208 3000
rect 105740 480 105768 2994
rect 106936 480 106964 2994
rect 108132 480 108160 2994
rect 109328 480 109356 2994
rect 111168 2854 111196 2994
rect 110512 2848 110564 2854
rect 110512 2790 110564 2796
rect 111156 2848 111208 2854
rect 111156 2790 111208 2796
rect 110524 480 110552 2790
rect 111628 480 111656 6886
rect 112824 480 112852 6886
rect 115124 2990 115152 6886
rect 115860 2990 115888 10270
rect 117240 2990 117268 326606
rect 119804 10396 119856 10402
rect 119804 10338 119856 10344
rect 119816 2990 119844 10338
rect 120000 6914 120028 328170
rect 119908 6886 120028 6914
rect 115112 2984 115164 2990
rect 115112 2926 115164 2932
rect 115204 2984 115256 2990
rect 115204 2926 115256 2932
rect 115848 2984 115900 2990
rect 115848 2926 115900 2932
rect 116400 2984 116452 2990
rect 116400 2926 116452 2932
rect 117228 2984 117280 2990
rect 117228 2926 117280 2932
rect 118792 2984 118844 2990
rect 118792 2926 118844 2932
rect 119804 2984 119856 2990
rect 119804 2926 119856 2932
rect 114008 2916 114060 2922
rect 114008 2858 114060 2864
rect 114020 480 114048 2858
rect 115216 480 115244 2926
rect 116412 480 116440 2926
rect 117596 2848 117648 2854
rect 117596 2790 117648 2796
rect 117608 480 117636 2790
rect 118804 480 118832 2926
rect 119908 480 119936 6886
rect 122116 2990 122144 337554
rect 124128 332308 124180 332314
rect 124128 332250 124180 332256
rect 122748 10464 122800 10470
rect 122748 10406 122800 10412
rect 122760 2990 122788 10406
rect 124140 2990 124168 332250
rect 125520 6914 125548 337622
rect 177302 336696 177358 336705
rect 177302 336631 177358 336640
rect 173162 336560 173218 336569
rect 173162 336495 173218 336504
rect 130382 336288 130438 336297
rect 130382 336223 130438 336232
rect 126888 335096 126940 335102
rect 126888 335038 126940 335044
rect 125428 6886 125548 6914
rect 125428 2990 125456 6886
rect 126900 2990 126928 335038
rect 129004 334824 129056 334830
rect 129004 334766 129056 334772
rect 128176 7676 128228 7682
rect 128176 7618 128228 7624
rect 122104 2984 122156 2990
rect 122104 2926 122156 2932
rect 122288 2984 122340 2990
rect 122288 2926 122340 2932
rect 122748 2984 122800 2990
rect 122748 2926 122800 2932
rect 123484 2984 123536 2990
rect 123484 2926 123536 2932
rect 124128 2984 124180 2990
rect 124128 2926 124180 2932
rect 124680 2984 124732 2990
rect 124680 2926 124732 2932
rect 125416 2984 125468 2990
rect 125416 2926 125468 2932
rect 125876 2984 125928 2990
rect 125876 2926 125928 2932
rect 126888 2984 126940 2990
rect 126888 2926 126940 2932
rect 126980 2984 127032 2990
rect 126980 2926 127032 2932
rect 121092 2916 121144 2922
rect 121092 2858 121144 2864
rect 121104 480 121132 2858
rect 122300 480 122328 2926
rect 123496 480 123524 2926
rect 124692 480 124720 2926
rect 125888 480 125916 2926
rect 126992 480 127020 2926
rect 128188 480 128216 7618
rect 129016 2990 129044 334766
rect 130396 6254 130424 336223
rect 151728 335300 151780 335306
rect 151728 335242 151780 335248
rect 147588 335232 147640 335238
rect 147588 335174 147640 335180
rect 144828 335164 144880 335170
rect 144828 335106 144880 335112
rect 140688 335028 140740 335034
rect 140688 334970 140740 334976
rect 137284 334960 137336 334966
rect 137284 334902 137336 334908
rect 133788 334892 133840 334898
rect 133788 334834 133840 334840
rect 131764 7744 131816 7750
rect 131764 7686 131816 7692
rect 130384 6248 130436 6254
rect 130384 6190 130436 6196
rect 130568 6248 130620 6254
rect 130568 6190 130620 6196
rect 129372 5092 129424 5098
rect 129372 5034 129424 5040
rect 129004 2984 129056 2990
rect 129004 2926 129056 2932
rect 129384 480 129412 5034
rect 130580 480 130608 6190
rect 131776 480 131804 7686
rect 133800 2854 133828 334834
rect 135168 333668 135220 333674
rect 135168 333610 135220 333616
rect 135180 2854 135208 333610
rect 135260 9172 135312 9178
rect 135260 9114 135312 9120
rect 132960 2848 133012 2854
rect 132960 2790 133012 2796
rect 133788 2848 133840 2854
rect 133788 2790 133840 2796
rect 134156 2848 134208 2854
rect 134156 2790 134208 2796
rect 135168 2848 135220 2854
rect 135168 2790 135220 2796
rect 132972 480 133000 2790
rect 134168 480 134196 2790
rect 135272 480 135300 9114
rect 137296 2854 137324 334902
rect 137928 332376 137980 332382
rect 137928 332318 137980 332324
rect 137940 6914 137968 332318
rect 138848 9240 138900 9246
rect 138848 9182 138900 9188
rect 137664 6886 137968 6914
rect 136456 2848 136508 2854
rect 136456 2790 136508 2796
rect 137284 2848 137336 2854
rect 137284 2790 137336 2796
rect 136468 480 136496 2790
rect 137664 480 137692 6886
rect 138860 480 138888 9182
rect 140700 2854 140728 334970
rect 144736 333736 144788 333742
rect 144736 333678 144788 333684
rect 142068 332444 142120 332450
rect 142068 332386 142120 332392
rect 142080 2854 142108 332386
rect 142436 9308 142488 9314
rect 142436 9250 142488 9256
rect 140044 2848 140096 2854
rect 140044 2790 140096 2796
rect 140688 2848 140740 2854
rect 140688 2790 140740 2796
rect 141240 2848 141292 2854
rect 141240 2790 141292 2796
rect 142068 2848 142120 2854
rect 142068 2790 142120 2796
rect 140056 480 140084 2790
rect 141252 480 141280 2790
rect 142448 480 142476 9250
rect 143540 2848 143592 2854
rect 143540 2790 143592 2796
rect 143552 480 143580 2790
rect 144748 480 144776 333678
rect 144840 2854 144868 335106
rect 146208 329724 146260 329730
rect 146208 329666 146260 329672
rect 146220 6914 146248 329666
rect 145944 6886 146248 6914
rect 144828 2848 144880 2854
rect 144828 2790 144880 2796
rect 145944 480 145972 6886
rect 147600 2854 147628 335174
rect 148968 332512 149020 332518
rect 148968 332454 149020 332460
rect 148980 2854 149008 332454
rect 150348 10532 150400 10538
rect 150348 10474 150400 10480
rect 150360 2854 150388 10474
rect 151740 2854 151768 335242
rect 155224 334552 155276 334558
rect 155224 334494 155276 334500
rect 153108 332580 153160 332586
rect 153108 332522 153160 332528
rect 153016 331152 153068 331158
rect 153016 331094 153068 331100
rect 147128 2848 147180 2854
rect 147128 2790 147180 2796
rect 147588 2848 147640 2854
rect 147588 2790 147640 2796
rect 148324 2848 148376 2854
rect 148324 2790 148376 2796
rect 148968 2848 149020 2854
rect 148968 2790 149020 2796
rect 149520 2848 149572 2854
rect 149520 2790 149572 2796
rect 150348 2848 150400 2854
rect 150348 2790 150400 2796
rect 150624 2848 150676 2854
rect 150624 2790 150676 2796
rect 151728 2848 151780 2854
rect 151728 2790 151780 2796
rect 151820 2848 151872 2854
rect 151820 2790 151872 2796
rect 147140 480 147168 2790
rect 148336 480 148364 2790
rect 149532 480 149560 2790
rect 150636 480 150664 2790
rect 151832 480 151860 2790
rect 153028 480 153056 331094
rect 153120 2854 153148 332522
rect 155236 2854 155264 334494
rect 158628 334484 158680 334490
rect 158628 334426 158680 334432
rect 155868 331832 155920 331838
rect 155868 331774 155920 331780
rect 155880 2854 155908 331774
rect 157248 17264 157300 17270
rect 157248 17206 157300 17212
rect 157260 2854 157288 17206
rect 158640 2854 158668 334426
rect 161388 334416 161440 334422
rect 161388 334358 161440 334364
rect 160100 9376 160152 9382
rect 160100 9318 160152 9324
rect 158904 7812 158956 7818
rect 158904 7754 158956 7760
rect 153108 2848 153160 2854
rect 153108 2790 153160 2796
rect 154212 2848 154264 2854
rect 154212 2790 154264 2796
rect 155224 2848 155276 2854
rect 155224 2790 155276 2796
rect 155408 2848 155460 2854
rect 155408 2790 155460 2796
rect 155868 2848 155920 2854
rect 155868 2790 155920 2796
rect 156604 2848 156656 2854
rect 156604 2790 156656 2796
rect 157248 2848 157300 2854
rect 157248 2790 157300 2796
rect 157800 2848 157852 2854
rect 157800 2790 157852 2796
rect 158628 2848 158680 2854
rect 158628 2790 158680 2796
rect 154224 480 154252 2790
rect 155420 480 155448 2790
rect 156616 480 156644 2790
rect 157812 480 157840 2790
rect 158916 480 158944 7754
rect 160112 480 160140 9318
rect 161400 6914 161428 334358
rect 169668 334348 169720 334354
rect 169668 334290 169720 334296
rect 166908 333872 166960 333878
rect 166908 333814 166960 333820
rect 162768 333804 162820 333810
rect 162768 333746 162820 333752
rect 162780 6914 162808 333746
rect 165528 11824 165580 11830
rect 165528 11766 165580 11772
rect 163688 7880 163740 7886
rect 163688 7822 163740 7828
rect 161308 6886 161428 6914
rect 162504 6886 162808 6914
rect 161308 480 161336 6886
rect 162504 480 162532 6886
rect 163700 480 163728 7822
rect 165540 2854 165568 11766
rect 166920 2854 166948 333814
rect 169576 333192 169628 333198
rect 169576 333134 169628 333140
rect 167184 7948 167236 7954
rect 167184 7890 167236 7896
rect 164884 2848 164936 2854
rect 164884 2790 164936 2796
rect 165528 2848 165580 2854
rect 165528 2790 165580 2796
rect 166080 2848 166132 2854
rect 166080 2790 166132 2796
rect 166908 2848 166960 2854
rect 166908 2790 166960 2796
rect 164896 480 164924 2790
rect 166092 480 166120 2790
rect 167196 480 167224 7890
rect 168380 2848 168432 2854
rect 168380 2790 168432 2796
rect 168392 480 168420 2790
rect 169588 480 169616 333134
rect 169680 2854 169708 334290
rect 173176 13122 173204 336495
rect 173164 13116 173216 13122
rect 173164 13058 173216 13064
rect 174268 8084 174320 8090
rect 174268 8026 174320 8032
rect 170772 8016 170824 8022
rect 170772 7958 170824 7964
rect 169668 2848 169720 2854
rect 169668 2790 169720 2796
rect 170784 480 170812 7958
rect 173164 6316 173216 6322
rect 173164 6258 173216 6264
rect 171968 5296 172020 5302
rect 171968 5238 172020 5244
rect 171980 480 172008 5238
rect 173176 480 173204 6258
rect 174280 480 174308 8026
rect 177316 7614 177344 336631
rect 180062 336424 180118 336433
rect 180062 336359 180118 336368
rect 206284 336388 206336 336394
rect 179328 332988 179380 332994
rect 179328 332930 179380 332936
rect 177304 7608 177356 7614
rect 177304 7550 177356 7556
rect 177856 7608 177908 7614
rect 177856 7550 177908 7556
rect 176660 6452 176712 6458
rect 176660 6394 176712 6400
rect 175464 5160 175516 5166
rect 175464 5102 175516 5108
rect 175476 480 175504 5102
rect 176672 480 176700 6394
rect 177868 480 177896 7550
rect 179340 6914 179368 332930
rect 179064 6886 179368 6914
rect 179064 480 179092 6886
rect 180076 6390 180104 336359
rect 206284 336330 206336 336336
rect 204904 336320 204956 336326
rect 204904 336262 204956 336268
rect 198004 336252 198056 336258
rect 198004 336194 198056 336200
rect 196624 336116 196676 336122
rect 196624 336058 196676 336064
rect 195244 336048 195296 336054
rect 195244 335990 195296 335996
rect 194416 334280 194468 334286
rect 194416 334222 194468 334228
rect 187608 333940 187660 333946
rect 187608 333882 187660 333888
rect 184848 331764 184900 331770
rect 184848 331706 184900 331712
rect 181444 8152 181496 8158
rect 181444 8094 181496 8100
rect 180064 6384 180116 6390
rect 180064 6326 180116 6332
rect 180248 6384 180300 6390
rect 180248 6326 180300 6332
rect 180260 480 180288 6326
rect 181456 480 181484 8094
rect 183744 6520 183796 6526
rect 183744 6462 183796 6468
rect 182548 5228 182600 5234
rect 182548 5170 182600 5176
rect 182560 480 182588 5170
rect 183756 480 183784 6462
rect 184860 3482 184888 331706
rect 187620 6914 187648 333882
rect 191748 333124 191800 333130
rect 191748 333066 191800 333072
rect 188988 331696 189040 331702
rect 188988 331638 189040 331644
rect 187344 6886 187648 6914
rect 186136 5364 186188 5370
rect 186136 5306 186188 5312
rect 184860 3454 184980 3482
rect 184952 480 184980 3454
rect 186148 480 186176 5306
rect 187344 480 187372 6886
rect 189000 2854 189028 331638
rect 189724 5432 189776 5438
rect 189724 5374 189776 5380
rect 188528 2848 188580 2854
rect 188528 2790 188580 2796
rect 188988 2848 189040 2854
rect 188988 2790 189040 2796
rect 188540 480 188568 2790
rect 189736 480 189764 5374
rect 191760 2854 191788 333066
rect 193128 331220 193180 331226
rect 193128 331162 193180 331168
rect 193140 2854 193168 331162
rect 193220 4208 193272 4214
rect 193220 4150 193272 4156
rect 190828 2848 190880 2854
rect 190828 2790 190880 2796
rect 191748 2848 191800 2854
rect 191748 2790 191800 2796
rect 192024 2848 192076 2854
rect 192024 2790 192076 2796
rect 193128 2848 193180 2854
rect 193128 2790 193180 2796
rect 190840 480 190868 2790
rect 192036 480 192064 2790
rect 193232 480 193260 4150
rect 194428 480 194456 334222
rect 195256 4214 195284 335990
rect 195888 330472 195940 330478
rect 195888 330414 195940 330420
rect 195900 6914 195928 330414
rect 195624 6886 195928 6914
rect 195244 4208 195296 4214
rect 195244 4150 195296 4156
rect 195624 480 195652 6886
rect 196636 5234 196664 336058
rect 196808 5568 196860 5574
rect 196808 5510 196860 5516
rect 196624 5228 196676 5234
rect 196624 5170 196676 5176
rect 196820 480 196848 5510
rect 198016 5166 198044 336194
rect 202144 336184 202196 336190
rect 202144 336126 202196 336132
rect 198648 333056 198700 333062
rect 198648 332998 198700 333004
rect 198004 5160 198056 5166
rect 198004 5102 198056 5108
rect 198660 2854 198688 332998
rect 199108 8220 199160 8226
rect 199108 8162 199160 8168
rect 197912 2848 197964 2854
rect 197912 2790 197964 2796
rect 198648 2848 198700 2854
rect 198648 2790 198700 2796
rect 197924 480 197952 2790
rect 199120 480 199148 8162
rect 201500 6588 201552 6594
rect 201500 6530 201552 6536
rect 200304 5160 200356 5166
rect 200304 5102 200356 5108
rect 200316 480 200344 5102
rect 201512 480 201540 6530
rect 202156 5574 202184 336126
rect 202788 330404 202840 330410
rect 202788 330346 202840 330352
rect 202800 6914 202828 330346
rect 202708 6886 202828 6914
rect 202144 5568 202196 5574
rect 202144 5510 202196 5516
rect 202708 480 202736 6886
rect 204916 5370 204944 336262
rect 205088 6656 205140 6662
rect 205088 6598 205140 6604
rect 204904 5364 204956 5370
rect 204904 5306 204956 5312
rect 203892 5228 203944 5234
rect 203892 5170 203944 5176
rect 203904 480 203932 5170
rect 205100 480 205128 6598
rect 206296 5302 206324 336330
rect 206928 332920 206980 332926
rect 206928 332862 206980 332868
rect 206284 5296 206336 5302
rect 206284 5238 206336 5244
rect 206940 2854 206968 332862
rect 209056 306338 209084 377062
rect 212448 334212 212500 334218
rect 212448 334154 212500 334160
rect 210976 332852 211028 332858
rect 210976 332794 211028 332800
rect 209044 306332 209096 306338
rect 209044 306274 209096 306280
rect 208584 6724 208636 6730
rect 208584 6666 208636 6672
rect 207388 5296 207440 5302
rect 207388 5238 207440 5244
rect 206192 2848 206244 2854
rect 206192 2790 206244 2796
rect 206928 2848 206980 2854
rect 206928 2790 206980 2796
rect 206204 480 206232 2790
rect 207400 480 207428 5238
rect 208596 480 208624 6666
rect 210988 2854 211016 332794
rect 212460 6914 212488 334154
rect 213196 45558 213224 378558
rect 214564 377188 214616 377194
rect 214564 377130 214616 377136
rect 213828 331628 213880 331634
rect 213828 331570 213880 331576
rect 213184 45552 213236 45558
rect 213184 45494 213236 45500
rect 212184 6886 212488 6914
rect 211068 5364 211120 5370
rect 211068 5306 211120 5312
rect 209780 2848 209832 2854
rect 209780 2790 209832 2796
rect 210976 2848 211028 2854
rect 210976 2790 211028 2796
rect 209792 480 209820 2790
rect 211080 2122 211108 5306
rect 210988 2094 211108 2122
rect 210988 480 211016 2094
rect 212184 480 212212 6886
rect 213840 2854 213868 331570
rect 214576 85542 214604 377130
rect 215956 189038 215984 378626
rect 220176 377392 220228 377398
rect 220176 377334 220228 377340
rect 220084 334144 220136 334150
rect 220084 334086 220136 334092
rect 216588 332784 216640 332790
rect 216588 332726 216640 332732
rect 215944 189032 215996 189038
rect 215944 188974 215996 188980
rect 214564 85536 214616 85542
rect 214564 85478 214616 85484
rect 215208 14476 215260 14482
rect 215208 14418 215260 14424
rect 215220 2854 215248 14418
rect 216600 2854 216628 332726
rect 217968 330336 218020 330342
rect 217968 330278 218020 330284
rect 217980 2854 218008 330278
rect 218060 5500 218112 5506
rect 218060 5442 218112 5448
rect 213368 2848 213420 2854
rect 213368 2790 213420 2796
rect 213828 2848 213880 2854
rect 213828 2790 213880 2796
rect 214472 2848 214524 2854
rect 214472 2790 214524 2796
rect 215208 2848 215260 2854
rect 215208 2790 215260 2796
rect 215668 2848 215720 2854
rect 215668 2790 215720 2796
rect 216588 2848 216640 2854
rect 216588 2790 216640 2796
rect 216864 2848 216916 2854
rect 216864 2790 216916 2796
rect 217968 2848 218020 2854
rect 217968 2790 218020 2796
rect 213380 480 213408 2790
rect 214484 480 214512 2790
rect 215680 480 215708 2790
rect 216876 480 216904 2790
rect 218072 480 218100 5442
rect 220096 2854 220124 334086
rect 220188 241466 220216 377334
rect 222844 336456 222896 336462
rect 222844 336398 222896 336404
rect 220728 330268 220780 330274
rect 220728 330210 220780 330216
rect 220176 241460 220228 241466
rect 220176 241402 220228 241408
rect 220740 6914 220768 330210
rect 222856 14482 222884 336398
rect 222948 293962 222976 379034
rect 228456 378956 228508 378962
rect 228456 378898 228508 378904
rect 224224 377732 224276 377738
rect 224224 377674 224276 377680
rect 224236 346390 224264 377674
rect 226984 377324 227036 377330
rect 226984 377266 227036 377272
rect 224224 346384 224276 346390
rect 224224 346326 224276 346332
rect 224224 336728 224276 336734
rect 224224 336670 224276 336676
rect 223488 332716 223540 332722
rect 223488 332658 223540 332664
rect 222936 293956 222988 293962
rect 222936 293898 222988 293904
rect 222844 14476 222896 14482
rect 222844 14418 222896 14424
rect 220464 6886 220768 6914
rect 219256 2848 219308 2854
rect 219256 2790 219308 2796
rect 220084 2848 220136 2854
rect 220084 2790 220136 2796
rect 219268 480 219296 2790
rect 220464 480 220492 6886
rect 221556 4752 221608 4758
rect 221556 4694 221608 4700
rect 221568 480 221596 4694
rect 223500 2854 223528 332658
rect 224236 11830 224264 336670
rect 224868 331560 224920 331566
rect 224868 331502 224920 331508
rect 224224 11824 224276 11830
rect 224224 11766 224276 11772
rect 224880 2854 224908 331502
rect 226996 33114 227024 377266
rect 228364 336524 228416 336530
rect 228364 336466 228416 336472
rect 227628 334076 227680 334082
rect 227628 334018 227680 334024
rect 227536 332648 227588 332654
rect 227536 332590 227588 332596
rect 226984 33108 227036 33114
rect 226984 33050 227036 33056
rect 227548 16574 227576 332590
rect 227456 16546 227576 16574
rect 225144 4208 225196 4214
rect 225144 4150 225196 4156
rect 222752 2848 222804 2854
rect 222752 2790 222804 2796
rect 223488 2848 223540 2854
rect 223488 2790 223540 2796
rect 223948 2848 224000 2854
rect 223948 2790 224000 2796
rect 224868 2848 224920 2854
rect 224868 2790 224920 2796
rect 222764 480 222792 2790
rect 223960 480 223988 2790
rect 225156 480 225184 4150
rect 227456 2854 227484 16546
rect 227640 6914 227668 334018
rect 227548 6886 227668 6914
rect 226340 2848 226392 2854
rect 226340 2790 226392 2796
rect 227444 2848 227496 2854
rect 227444 2790 227496 2796
rect 226352 480 226380 2790
rect 227548 480 227576 6886
rect 228376 4214 228404 336466
rect 228468 71738 228496 378898
rect 231124 335912 231176 335918
rect 231124 335854 231176 335860
rect 230480 335572 230532 335578
rect 230480 335514 230532 335520
rect 230492 334354 230520 335514
rect 230480 334348 230532 334354
rect 230480 334290 230532 334296
rect 230388 334008 230440 334014
rect 230388 333950 230440 333956
rect 228456 71732 228508 71738
rect 228456 71674 228508 71680
rect 228732 13116 228784 13122
rect 228732 13058 228784 13064
rect 228364 4208 228416 4214
rect 228364 4150 228416 4156
rect 228744 480 228772 13058
rect 230400 3534 230428 333950
rect 231032 9444 231084 9450
rect 231032 9386 231084 9392
rect 229836 3528 229888 3534
rect 229836 3470 229888 3476
rect 230388 3528 230440 3534
rect 230388 3470 230440 3476
rect 229848 480 229876 3470
rect 231044 480 231072 9386
rect 231136 4758 231164 335854
rect 231228 215286 231256 379170
rect 231768 335980 231820 335986
rect 231768 335922 231820 335928
rect 231676 335368 231728 335374
rect 231676 335310 231728 335316
rect 231216 215280 231268 215286
rect 231216 215222 231268 215228
rect 231124 4752 231176 4758
rect 231124 4694 231176 4700
rect 231688 4690 231716 335310
rect 231676 4684 231728 4690
rect 231676 4626 231728 4632
rect 231780 4554 231808 335922
rect 232504 335844 232556 335850
rect 232504 335786 232556 335792
rect 232516 5506 232544 335786
rect 232608 267714 232636 379238
rect 233056 336592 233108 336598
rect 233056 336534 233108 336540
rect 232596 267708 232648 267714
rect 232596 267650 232648 267656
rect 233068 5506 233096 336534
rect 233976 335776 234028 335782
rect 233976 335718 234028 335724
rect 233884 335708 233936 335714
rect 233884 335650 233936 335656
rect 233148 335504 233200 335510
rect 233148 335446 233200 335452
rect 233160 334422 233188 335446
rect 233424 335436 233476 335442
rect 233424 335378 233476 335384
rect 233148 334416 233200 334422
rect 233148 334358 233200 334364
rect 233240 334348 233292 334354
rect 233240 334290 233292 334296
rect 233252 334234 233280 334290
rect 233160 334206 233280 334234
rect 232504 5500 232556 5506
rect 232504 5442 232556 5448
rect 233056 5500 233108 5506
rect 233056 5442 233108 5448
rect 231768 4548 231820 4554
rect 231768 4490 231820 4496
rect 233160 3534 233188 334206
rect 233436 332994 233464 335378
rect 233424 332988 233476 332994
rect 233424 332930 233476 332936
rect 233896 5438 233924 335650
rect 233988 13122 234016 335718
rect 234080 320142 234108 379374
rect 243360 379364 243412 379370
rect 243360 379306 243412 379312
rect 242348 379024 242400 379030
rect 242348 378966 242400 378972
rect 239680 378412 239732 378418
rect 239680 378354 239732 378360
rect 237196 378276 237248 378282
rect 237196 378218 237248 378224
rect 237104 378208 237156 378214
rect 237104 378150 237156 378156
rect 237116 377890 237144 378150
rect 236808 377862 237144 377890
rect 237208 377754 237236 378218
rect 239692 377890 239720 378354
rect 240048 378344 240100 378350
rect 240048 378286 240100 378292
rect 240060 377890 240088 378286
rect 242360 377890 242388 378966
rect 243372 377890 243400 379306
rect 248052 379160 248104 379166
rect 248052 379102 248104 379108
rect 245476 378888 245528 378894
rect 245476 378830 245528 378836
rect 244924 377936 244976 377942
rect 239384 377862 239720 377890
rect 239936 377862 240088 377890
rect 242052 377862 242388 377890
rect 243064 377862 243400 377890
rect 244628 377884 244924 377890
rect 245488 377890 245516 378830
rect 246028 378820 246080 378826
rect 246028 378762 246080 378768
rect 246040 377890 246068 378762
rect 248064 377890 248092 379102
rect 249156 378752 249208 378758
rect 249156 378694 249208 378700
rect 248236 378480 248288 378486
rect 248236 378422 248288 378428
rect 244628 377878 244976 377884
rect 244628 377862 244964 377878
rect 245180 377862 245516 377890
rect 245732 377862 246068 377890
rect 246284 377874 246620 377890
rect 246284 377868 246632 377874
rect 246284 377862 246580 377868
rect 247848 377862 248092 377890
rect 248248 377890 248276 378422
rect 249168 377890 249196 378694
rect 249720 377890 249748 404330
rect 250916 383654 250944 418134
rect 250824 383626 250944 383654
rect 250260 379704 250312 379710
rect 250260 379646 250312 379652
rect 250272 377890 250300 379646
rect 250824 377890 250852 383626
rect 251008 379710 251036 430578
rect 250996 379704 251048 379710
rect 250996 379646 251048 379652
rect 251100 377890 251128 456758
rect 251824 379704 251876 379710
rect 251824 379646 251876 379652
rect 251836 377890 251864 379646
rect 252296 377890 252324 470562
rect 252388 379710 252416 484366
rect 252376 379704 252428 379710
rect 252376 379646 252428 379652
rect 248248 377862 248308 377890
rect 248860 377862 249196 377890
rect 249412 377862 249748 377890
rect 249964 377862 250300 377890
rect 250424 377862 250852 377890
rect 250976 377862 251128 377890
rect 251528 377862 251864 377890
rect 252080 377862 252324 377890
rect 252480 377890 252508 510614
rect 253388 379704 253440 379710
rect 253388 379646 253440 379652
rect 253400 377890 253428 379646
rect 253768 377890 253796 524418
rect 253860 379710 253888 536794
rect 255056 379710 255084 563042
rect 253848 379704 253900 379710
rect 253848 379646 253900 379652
rect 254400 379704 254452 379710
rect 254400 379646 254452 379652
rect 255044 379704 255096 379710
rect 255044 379646 255096 379652
rect 254412 377890 254440 379646
rect 254952 379568 255004 379574
rect 254952 379510 255004 379516
rect 254964 377890 254992 379510
rect 252480 377862 252540 377890
rect 253092 377862 253428 377890
rect 253644 377862 253796 377890
rect 254104 377862 254440 377890
rect 254656 377862 254992 377890
rect 255148 377890 255176 576846
rect 255240 379574 255268 590650
rect 256528 379710 256556 616830
rect 256056 379704 256108 379710
rect 256056 379646 256108 379652
rect 256516 379704 256568 379710
rect 256516 379646 256568 379652
rect 255228 379568 255280 379574
rect 255228 379510 255280 379516
rect 256068 377890 256096 379646
rect 256620 377890 256648 643078
rect 257804 630692 257856 630698
rect 257804 630634 257856 630640
rect 257816 379710 257844 630634
rect 257068 379704 257120 379710
rect 257068 379646 257120 379652
rect 257804 379704 257856 379710
rect 257804 379646 257856 379652
rect 257080 377890 257108 379646
rect 257908 378162 257936 670686
rect 257632 378134 257936 378162
rect 257632 377890 257660 378134
rect 258000 377890 258028 696934
rect 259184 683188 259236 683194
rect 259184 683130 259236 683136
rect 259196 379846 259224 683130
rect 258632 379840 258684 379846
rect 258632 379782 258684 379788
rect 259184 379840 259236 379846
rect 259184 379782 259236 379788
rect 258644 377890 258672 379782
rect 259288 377890 259316 700266
rect 255148 377862 255208 377890
rect 255760 377862 256096 377890
rect 256220 377862 256648 377890
rect 256772 377862 257108 377890
rect 257324 377862 257660 377890
rect 257784 377862 258028 377890
rect 258336 377862 258672 377890
rect 258888 377862 259316 377890
rect 259380 377890 259408 700402
rect 260196 379840 260248 379846
rect 260196 379782 260248 379788
rect 260208 377890 260236 379782
rect 260668 377890 260696 700538
rect 260748 700392 260800 700398
rect 260748 700334 260800 700340
rect 260760 379846 260788 700334
rect 261956 383654 261984 700606
rect 261864 383626 261984 383654
rect 260748 379840 260800 379846
rect 260748 379782 260800 379788
rect 261300 379840 261352 379846
rect 261300 379782 261352 379788
rect 261312 377890 261340 379782
rect 261864 377890 261892 383626
rect 262048 378162 262076 700810
rect 262128 700732 262180 700738
rect 262128 700674 262180 700680
rect 262140 379846 262168 700674
rect 263336 379846 263364 700946
rect 263508 700936 263560 700942
rect 263508 700878 263560 700884
rect 263416 700188 263468 700194
rect 263416 700130 263468 700136
rect 262128 379840 262180 379846
rect 262128 379782 262180 379788
rect 262864 379840 262916 379846
rect 262864 379782 262916 379788
rect 263324 379840 263376 379846
rect 263324 379782 263376 379788
rect 259380 377862 259440 377890
rect 259900 377862 260236 377890
rect 260452 377862 260696 377890
rect 261004 377862 261340 377890
rect 261464 377862 261892 377890
rect 262002 378134 262076 378162
rect 262002 377876 262030 378134
rect 262876 377890 262904 379782
rect 263324 379636 263376 379642
rect 263324 379578 263376 379584
rect 263336 377890 263364 379578
rect 262568 377862 262904 377890
rect 263120 377862 263364 377890
rect 263428 377890 263456 700130
rect 263520 379642 263548 700878
rect 264796 700120 264848 700126
rect 264796 700062 264848 700068
rect 264428 379704 264480 379710
rect 264428 379646 264480 379652
rect 263508 379636 263560 379642
rect 263508 379578 263560 379584
rect 264440 377890 264468 379646
rect 264808 377890 264836 700062
rect 264888 700052 264940 700058
rect 264888 699994 264940 700000
rect 264900 379710 264928 699994
rect 266452 699984 266504 699990
rect 266452 699926 266504 699932
rect 266268 699712 266320 699718
rect 266268 699654 266320 699660
rect 266280 383654 266308 699654
rect 266464 402974 266492 699926
rect 267660 699718 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 269488 700800 269540 700806
rect 269488 700742 269540 700748
rect 267924 700256 267976 700262
rect 267924 700198 267976 700204
rect 267648 699712 267700 699718
rect 267648 699654 267700 699660
rect 267936 402974 267964 700198
rect 269500 402974 269528 700742
rect 271880 700528 271932 700534
rect 271880 700470 271932 700476
rect 266464 402946 266952 402974
rect 267936 402946 268516 402974
rect 269500 402946 270080 402974
rect 266096 383626 266308 383654
rect 264888 379704 264940 379710
rect 264888 379646 264940 379652
rect 265532 379704 265584 379710
rect 265532 379646 265584 379652
rect 265544 377890 265572 379646
rect 266096 377890 266124 383626
rect 266452 379636 266504 379642
rect 266452 379578 266504 379584
rect 266268 379568 266320 379574
rect 266268 379510 266320 379516
rect 266280 378162 266308 379510
rect 263428 377862 263580 377890
rect 264132 377862 264468 377890
rect 264684 377862 264836 377890
rect 265236 377862 265572 377890
rect 265696 377862 266124 377890
rect 266188 378134 266308 378162
rect 246580 377810 246632 377816
rect 243912 377800 243964 377806
rect 237208 377726 237268 377754
rect 243616 377748 243912 377754
rect 243616 377742 243964 377748
rect 266188 377754 266216 378134
rect 266464 377890 266492 379578
rect 266924 377890 266952 402946
rect 267740 379840 267792 379846
rect 267740 379782 267792 379788
rect 267752 377890 267780 379782
rect 268016 379772 268068 379778
rect 268016 379714 268068 379720
rect 268028 377890 268056 379714
rect 268488 377890 268516 402946
rect 269580 380044 269632 380050
rect 269580 379986 269632 379992
rect 269120 379908 269172 379914
rect 269120 379850 269172 379856
rect 269132 377890 269160 379850
rect 269592 377890 269620 379986
rect 270052 377890 270080 402946
rect 271144 380112 271196 380118
rect 271144 380054 271196 380060
rect 270592 379976 270644 379982
rect 270592 379918 270644 379924
rect 270604 377890 270632 379918
rect 271156 377890 271184 380054
rect 271788 379636 271840 379642
rect 271788 379578 271840 379584
rect 266464 377862 266800 377890
rect 266924 377862 267260 377890
rect 267752 377862 267812 377890
rect 268028 377862 268364 377890
rect 268488 377862 268916 377890
rect 269132 377862 269376 377890
rect 269592 377862 269928 377890
rect 270052 377862 270480 377890
rect 270604 377862 270940 377890
rect 271156 377862 271492 377890
rect 243616 377726 243952 377742
rect 266188 377726 266248 377754
rect 246948 377664 247000 377670
rect 238372 377602 238616 377618
rect 238924 377602 239260 377618
rect 240488 377602 240824 377618
rect 241500 377602 241652 377618
rect 246744 377612 246948 377618
rect 246744 377606 247000 377612
rect 238372 377596 238628 377602
rect 238372 377590 238576 377596
rect 238924 377596 239272 377602
rect 238924 377590 239220 377596
rect 238576 377538 238628 377544
rect 240488 377596 240836 377602
rect 240488 377590 240784 377596
rect 239220 377538 239272 377544
rect 241500 377596 241664 377602
rect 241500 377590 241612 377596
rect 240784 377538 240836 377544
rect 246744 377590 246988 377606
rect 247296 377602 247632 377618
rect 247296 377596 247644 377602
rect 247296 377590 247592 377596
rect 241612 377538 241664 377544
rect 247592 377538 247644 377544
rect 271800 377534 271828 379578
rect 271892 377890 271920 700470
rect 273444 656940 273496 656946
rect 273444 656882 273496 656888
rect 272246 380352 272302 380361
rect 272246 380287 272302 380296
rect 272260 377890 272288 380287
rect 272706 380216 272762 380225
rect 272706 380151 272762 380160
rect 272720 377890 272748 380151
rect 273456 377890 273484 656882
rect 274732 605872 274784 605878
rect 274732 605814 274784 605820
rect 274272 380860 274324 380866
rect 274272 380802 274324 380808
rect 273812 380792 273864 380798
rect 273812 380734 273864 380740
rect 273824 377890 273852 380734
rect 274284 377890 274312 380802
rect 274744 377890 274772 605814
rect 276388 553444 276440 553450
rect 276388 553386 276440 553392
rect 275376 380724 275428 380730
rect 275376 380666 275428 380672
rect 275388 377890 275416 380666
rect 276020 380588 276072 380594
rect 276020 380530 276072 380536
rect 276032 377890 276060 380530
rect 276400 377890 276428 553386
rect 277492 501016 277544 501022
rect 277492 500958 277544 500964
rect 277504 402974 277532 500958
rect 278964 448588 279016 448594
rect 278964 448530 279016 448536
rect 278976 402974 279004 448530
rect 277504 402946 277992 402974
rect 278976 402946 279556 402974
rect 276940 380656 276992 380662
rect 276940 380598 276992 380604
rect 276952 377890 276980 380598
rect 277584 380520 277636 380526
rect 277584 380462 277636 380468
rect 277596 377890 277624 380462
rect 277964 377890 277992 402946
rect 278780 380452 278832 380458
rect 278780 380394 278832 380400
rect 278792 377890 278820 380394
rect 279056 380384 279108 380390
rect 279056 380326 279108 380332
rect 279068 377890 279096 380326
rect 279528 377890 279556 402946
rect 281080 397520 281132 397526
rect 281080 397462 281132 397468
rect 280160 380316 280212 380322
rect 280160 380258 280212 380264
rect 280172 377890 280200 380258
rect 280620 380248 280672 380254
rect 280620 380190 280672 380196
rect 280528 379772 280580 379778
rect 280528 379714 280580 379720
rect 271892 377862 272044 377890
rect 272260 377862 272596 377890
rect 272720 377862 273056 377890
rect 273456 377862 273608 377890
rect 273824 377862 274160 377890
rect 274284 377862 274620 377890
rect 274744 377862 275172 377890
rect 275388 377862 275724 377890
rect 276032 377862 276276 377890
rect 276400 377862 276736 377890
rect 276952 377862 277288 377890
rect 277596 377862 277840 377890
rect 277964 377862 278300 377890
rect 278792 377862 278852 377890
rect 279068 377862 279404 377890
rect 279528 377862 279956 377890
rect 280172 377862 280416 377890
rect 271788 377528 271840 377534
rect 271788 377470 271840 377476
rect 280540 377466 280568 379714
rect 280632 377890 280660 380190
rect 281092 377890 281120 397462
rect 281724 380180 281776 380186
rect 281724 380122 281776 380128
rect 281736 377890 281764 380122
rect 282932 379574 282960 702406
rect 290096 379772 290148 379778
rect 290096 379714 290148 379720
rect 283288 379636 283340 379642
rect 283288 379578 283340 379584
rect 282920 379568 282972 379574
rect 282920 379510 282972 379516
rect 282184 378548 282236 378554
rect 282184 378490 282236 378496
rect 282196 377890 282224 378490
rect 283300 377890 283328 379578
rect 283748 379432 283800 379438
rect 283748 379374 283800 379380
rect 283760 377890 283788 379374
rect 285680 379296 285732 379302
rect 285680 379238 285732 379244
rect 284300 379092 284352 379098
rect 284300 379034 284352 379040
rect 284312 377890 284340 379034
rect 285692 377890 285720 379238
rect 287152 379228 287204 379234
rect 287152 379170 287204 379176
rect 287164 377890 287192 379170
rect 287428 378684 287480 378690
rect 287428 378626 287480 378632
rect 287440 377890 287468 378626
rect 290108 377890 290136 379714
rect 299492 379710 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 700058 332548 703520
rect 348804 700126 348832 703520
rect 364996 700194 365024 703520
rect 397472 701010 397500 703520
rect 397460 701004 397512 701010
rect 397460 700946 397512 700952
rect 413664 700942 413692 703520
rect 413652 700936 413704 700942
rect 413652 700878 413704 700884
rect 429856 700874 429884 703520
rect 429844 700868 429896 700874
rect 429844 700810 429896 700816
rect 462332 700738 462360 703520
rect 462320 700732 462372 700738
rect 462320 700674 462372 700680
rect 478524 700670 478552 703520
rect 478512 700664 478564 700670
rect 478512 700606 478564 700612
rect 494808 700602 494836 703520
rect 494796 700596 494848 700602
rect 494796 700538 494848 700544
rect 527192 700466 527220 703520
rect 527180 700460 527232 700466
rect 527180 700402 527232 700408
rect 543476 700398 543504 703520
rect 543464 700392 543516 700398
rect 543464 700334 543516 700340
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 364984 700188 365036 700194
rect 364984 700130 365036 700136
rect 348792 700120 348844 700126
rect 348792 700062 348844 700068
rect 332508 700052 332560 700058
rect 332508 699994 332560 700000
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 299480 379704 299532 379710
rect 299480 379646 299532 379652
rect 295984 379364 296036 379370
rect 295984 379306 296036 379312
rect 291660 378956 291712 378962
rect 291660 378898 291712 378904
rect 291672 377890 291700 378898
rect 292212 378616 292264 378622
rect 292212 378558 292264 378564
rect 292224 377890 292252 378558
rect 280632 377862 280968 377890
rect 281092 377862 281520 377890
rect 281736 377862 282072 377890
rect 282196 377862 282532 377890
rect 283300 377862 283636 377890
rect 283760 377862 284096 377890
rect 284312 377862 284648 377890
rect 285692 377862 285752 377890
rect 287164 377862 287316 377890
rect 287440 377862 287776 377890
rect 290108 377862 290444 377890
rect 291672 377862 292008 377890
rect 292224 377862 292560 377890
rect 282932 377738 283084 377754
rect 282920 377732 283084 377738
rect 282972 377726 283084 377732
rect 282920 377674 282972 377680
rect 284864 377466 285200 377482
rect 280528 377460 280580 377466
rect 280528 377402 280580 377408
rect 284852 377460 285200 377466
rect 284904 377454 285200 377460
rect 284852 377402 284904 377408
rect 285864 377392 285916 377398
rect 235446 377360 235502 377369
rect 234632 377318 235244 377346
rect 234526 335880 234582 335889
rect 234526 335815 234582 335824
rect 234436 335640 234488 335646
rect 234436 335582 234488 335588
rect 234344 331492 234396 331498
rect 234344 331434 234396 331440
rect 234356 325694 234384 331434
rect 234448 330562 234476 335582
rect 234540 335102 234568 335815
rect 234528 335096 234580 335102
rect 234528 335038 234580 335044
rect 234448 330534 234568 330562
rect 234356 325666 234476 325694
rect 234068 320136 234120 320142
rect 234068 320078 234120 320084
rect 233976 13116 234028 13122
rect 233976 13058 234028 13064
rect 233884 5432 233936 5438
rect 233884 5374 233936 5380
rect 234448 3534 234476 325666
rect 234540 4214 234568 330534
rect 234632 6866 234660 377318
rect 236550 377360 236606 377369
rect 235502 377318 235704 377346
rect 236256 377318 236550 377346
rect 235446 377295 235502 377304
rect 238114 377360 238170 377369
rect 237820 377318 238114 377346
rect 236550 377295 236606 377304
rect 241242 377360 241298 377369
rect 240948 377318 241242 377346
rect 238114 377295 238170 377304
rect 242714 377360 242770 377369
rect 242604 377318 242714 377346
rect 241242 377295 241298 377304
rect 242714 377295 242770 377304
rect 244002 377360 244058 377369
rect 244058 377318 244168 377346
rect 288532 377392 288584 377398
rect 286414 377360 286470 377369
rect 285916 377340 286212 377346
rect 285864 377334 286212 377340
rect 285876 377318 286212 377334
rect 244002 377295 244058 377304
rect 287978 377360 288034 377369
rect 286470 377318 286764 377346
rect 286414 377295 286470 377304
rect 288034 377318 288328 377346
rect 290648 377392 290700 377398
rect 289082 377360 289138 377369
rect 288584 377340 288880 377346
rect 288532 377334 288880 377340
rect 288544 377318 288880 377334
rect 287978 377295 288034 377304
rect 290186 377360 290242 377369
rect 289138 377318 289432 377346
rect 289892 377318 290186 377346
rect 289082 377295 289138 377304
rect 293224 377392 293276 377398
rect 291198 377360 291254 377369
rect 290700 377340 290996 377346
rect 290648 377334 290996 377340
rect 290660 377318 290996 377334
rect 290186 377295 290242 377304
rect 292762 377360 292818 377369
rect 291254 377318 291456 377346
rect 291198 377295 291254 377304
rect 292818 377318 293112 377346
rect 294326 377360 294382 377369
rect 293276 377340 293572 377346
rect 293224 377334 293572 377340
rect 293236 377318 293572 377334
rect 294124 377318 294326 377346
rect 292762 377295 292818 377304
rect 294676 377318 295104 377346
rect 294326 377295 294382 377304
rect 234710 377224 234766 377233
rect 234710 377159 234766 377168
rect 294970 377224 295026 377233
rect 294970 377159 295026 377168
rect 234724 33114 234752 377159
rect 294984 340874 295012 377159
rect 295076 345014 295104 377318
rect 295076 344986 295288 345014
rect 294984 340846 295196 340874
rect 235000 338014 235060 338042
rect 234804 337884 234856 337890
rect 234804 337826 234856 337832
rect 234712 33108 234764 33114
rect 234712 33050 234764 33056
rect 234620 6860 234672 6866
rect 234620 6802 234672 6808
rect 234620 5024 234672 5030
rect 234620 4966 234672 4972
rect 234528 4208 234580 4214
rect 234528 4150 234580 4156
rect 232228 3528 232280 3534
rect 232228 3470 232280 3476
rect 233148 3528 233200 3534
rect 233148 3470 233200 3476
rect 233424 3528 233476 3534
rect 233424 3470 233476 3476
rect 234436 3528 234488 3534
rect 234436 3470 234488 3476
rect 232240 480 232268 3470
rect 233436 480 233464 3470
rect 234632 480 234660 4966
rect 234816 3369 234844 337826
rect 235000 326738 235028 338014
rect 235138 337770 235166 338028
rect 235092 337742 235166 337770
rect 234988 326732 235040 326738
rect 234988 326674 235040 326680
rect 235092 326448 235120 337742
rect 235230 337634 235258 338028
rect 235322 337770 235350 338028
rect 235460 338014 235520 338042
rect 235322 337742 235396 337770
rect 234908 326420 235120 326448
rect 235184 337606 235258 337634
rect 234908 4894 234936 326420
rect 235184 326346 235212 337606
rect 235368 328454 235396 337742
rect 235460 336569 235488 338014
rect 235598 337890 235626 338028
rect 235586 337884 235638 337890
rect 235586 337826 235638 337832
rect 235690 337770 235718 338028
rect 235644 337742 235718 337770
rect 235828 338014 235888 338042
rect 235446 336560 235502 336569
rect 235446 336495 235502 336504
rect 235092 326318 235212 326346
rect 235276 328426 235396 328454
rect 234988 323604 235040 323610
rect 234988 323546 235040 323552
rect 234896 4888 234948 4894
rect 234896 4830 234948 4836
rect 235000 4758 235028 323546
rect 235092 4826 235120 326318
rect 235172 326256 235224 326262
rect 235172 326198 235224 326204
rect 235184 4962 235212 326198
rect 235276 6186 235304 328426
rect 235644 326262 235672 337742
rect 235632 326256 235684 326262
rect 235632 326198 235684 326204
rect 235828 316034 235856 338014
rect 235966 337770 235994 338028
rect 236058 337906 236086 338028
rect 236196 338014 236256 338042
rect 236058 337878 236132 337906
rect 235920 337742 235994 337770
rect 235920 336705 235948 337742
rect 235906 336696 235962 336705
rect 235906 336631 235962 336640
rect 236104 336025 236132 337878
rect 236196 336802 236224 338014
rect 236334 337770 236362 338028
rect 236288 337742 236362 337770
rect 236184 336796 236236 336802
rect 236184 336738 236236 336744
rect 236090 336016 236146 336025
rect 236090 335951 236146 335960
rect 236288 330614 236316 337742
rect 236426 337668 236454 338028
rect 236380 337640 236454 337668
rect 236564 338014 236624 338042
rect 236276 330608 236328 330614
rect 236276 330550 236328 330556
rect 236184 326392 236236 326398
rect 236184 326334 236236 326340
rect 235368 316006 235856 316034
rect 235368 8974 235396 316006
rect 235356 8968 235408 8974
rect 235356 8910 235408 8916
rect 235264 6180 235316 6186
rect 235264 6122 235316 6128
rect 235172 4956 235224 4962
rect 235172 4898 235224 4904
rect 235080 4820 235132 4826
rect 235080 4762 235132 4768
rect 234988 4752 235040 4758
rect 234988 4694 235040 4700
rect 235816 4208 235868 4214
rect 235816 4150 235868 4156
rect 234802 3360 234858 3369
rect 234802 3295 234858 3304
rect 235828 480 235856 4150
rect 236196 3641 236224 326334
rect 236182 3632 236238 3641
rect 236182 3567 236238 3576
rect 236380 3505 236408 337640
rect 236564 326398 236592 338014
rect 236702 337770 236730 338028
rect 236794 337906 236822 338028
rect 236932 338014 236992 338042
rect 236794 337878 236868 337906
rect 236656 337742 236730 337770
rect 236656 334626 236684 337742
rect 236644 334620 236696 334626
rect 236644 334562 236696 334568
rect 236840 329186 236868 337878
rect 236932 336161 236960 338014
rect 237070 337770 237098 338028
rect 237162 337906 237190 338028
rect 237300 338014 237360 338042
rect 237162 337878 237236 337906
rect 237024 337742 237098 337770
rect 236918 336152 236974 336161
rect 236918 336087 236974 336096
rect 236828 329180 236880 329186
rect 236828 329122 236880 329128
rect 236552 326392 236604 326398
rect 236552 326334 236604 326340
rect 237024 316034 237052 337742
rect 237208 333266 237236 337878
rect 237196 333260 237248 333266
rect 237196 333202 237248 333208
rect 237300 327894 237328 338014
rect 237438 337770 237466 338028
rect 237392 337742 237466 337770
rect 237530 337770 237558 338028
rect 237668 338014 237728 338042
rect 237530 337742 237604 337770
rect 237288 327888 237340 327894
rect 237288 327830 237340 327836
rect 237392 326398 237420 337742
rect 237472 334620 237524 334626
rect 237472 334562 237524 334568
rect 237484 327758 237512 334562
rect 237576 328454 237604 337742
rect 237668 336870 237696 338014
rect 237806 337906 237834 338028
rect 237760 337878 237834 337906
rect 237656 336864 237708 336870
rect 237656 336806 237708 336812
rect 237760 334626 237788 337878
rect 237898 337770 237926 338028
rect 237852 337742 237926 337770
rect 238036 338014 238096 338042
rect 237852 336297 237880 337742
rect 237932 337680 237984 337686
rect 237932 337622 237984 337628
rect 237838 336288 237894 336297
rect 237838 336223 237894 336232
rect 237748 334620 237800 334626
rect 237748 334562 237800 334568
rect 237944 331214 237972 337622
rect 238036 331974 238064 338014
rect 238174 337770 238202 338028
rect 238128 337742 238202 337770
rect 238024 331968 238076 331974
rect 238024 331910 238076 331916
rect 237852 331186 237972 331214
rect 237576 328426 237696 328454
rect 237472 327752 237524 327758
rect 237472 327694 237524 327700
rect 237380 326392 237432 326398
rect 237380 326334 237432 326340
rect 236564 316006 237052 316034
rect 236564 3777 236592 316006
rect 237012 4820 237064 4826
rect 237012 4762 237064 4768
rect 236550 3768 236606 3777
rect 236550 3703 236606 3712
rect 236366 3496 236422 3505
rect 236366 3431 236422 3440
rect 237024 480 237052 4762
rect 237668 3466 237696 328426
rect 237852 3602 237880 331186
rect 238128 329118 238156 337742
rect 238266 337668 238294 338028
rect 238220 337640 238294 337668
rect 238404 338014 238464 338042
rect 238116 329112 238168 329118
rect 238116 329054 238168 329060
rect 237932 326392 237984 326398
rect 237932 326334 237984 326340
rect 237840 3596 237892 3602
rect 237840 3538 237892 3544
rect 237656 3460 237708 3466
rect 237656 3402 237708 3408
rect 237944 2854 237972 326334
rect 238220 316034 238248 337640
rect 238404 336938 238432 338014
rect 238542 337770 238570 338028
rect 238634 337890 238662 338028
rect 238622 337884 238674 337890
rect 238622 337826 238674 337832
rect 238726 337770 238754 338028
rect 238496 337742 238570 337770
rect 238680 337742 238754 337770
rect 238910 337770 238938 338028
rect 239002 337958 239030 338028
rect 238990 337952 239042 337958
rect 238990 337894 239042 337900
rect 239094 337906 239122 338028
rect 239094 337878 239168 337906
rect 239036 337816 239088 337822
rect 238910 337742 238984 337770
rect 239036 337758 239088 337764
rect 238392 336932 238444 336938
rect 238392 336874 238444 336880
rect 238496 326466 238524 337742
rect 238680 331214 238708 337742
rect 238588 331186 238708 331214
rect 238588 330206 238616 331186
rect 238956 330682 238984 337742
rect 238944 330676 238996 330682
rect 238944 330618 238996 330624
rect 238576 330200 238628 330206
rect 238576 330142 238628 330148
rect 238484 326460 238536 326466
rect 238484 326402 238536 326408
rect 239048 326398 239076 337758
rect 239140 337006 239168 337878
rect 239278 337770 239306 338028
rect 239370 337958 239398 338028
rect 239358 337952 239410 337958
rect 239358 337894 239410 337900
rect 239462 337872 239490 338028
rect 239600 338014 239660 338042
rect 239462 337844 239536 337872
rect 239278 337742 239352 337770
rect 239220 337680 239272 337686
rect 239220 337622 239272 337628
rect 239128 337000 239180 337006
rect 239128 336942 239180 336948
rect 239128 334620 239180 334626
rect 239128 334562 239180 334568
rect 239036 326392 239088 326398
rect 239036 326334 239088 326340
rect 238128 316006 238248 316034
rect 238128 6914 238156 316006
rect 238036 6886 238156 6914
rect 238036 3806 238064 6886
rect 238116 4956 238168 4962
rect 238116 4898 238168 4904
rect 238024 3800 238076 3806
rect 238024 3742 238076 3748
rect 237932 2848 237984 2854
rect 237932 2790 237984 2796
rect 238128 480 238156 4898
rect 239140 3874 239168 334562
rect 239128 3868 239180 3874
rect 239128 3810 239180 3816
rect 239232 3738 239260 337622
rect 239324 333538 239352 337742
rect 239508 337142 239536 337844
rect 239496 337136 239548 337142
rect 239496 337078 239548 337084
rect 239312 333532 239364 333538
rect 239312 333474 239364 333480
rect 239600 331214 239628 338014
rect 239738 337770 239766 338028
rect 239830 337906 239858 338028
rect 239968 338014 240028 338042
rect 239830 337878 239904 337906
rect 239692 337742 239766 337770
rect 239692 334626 239720 337742
rect 239876 337074 239904 337878
rect 239864 337068 239916 337074
rect 239864 337010 239916 337016
rect 239680 334620 239732 334626
rect 239680 334562 239732 334568
rect 239968 332042 239996 338014
rect 240106 337770 240134 338028
rect 240198 337906 240226 338028
rect 240336 338014 240396 338042
rect 240198 337878 240272 337906
rect 240060 337742 240134 337770
rect 239956 332036 240008 332042
rect 239956 331978 240008 331984
rect 239324 331186 239628 331214
rect 239324 327826 239352 331186
rect 239312 327820 239364 327826
rect 239312 327762 239364 327768
rect 240060 326534 240088 337742
rect 240244 334694 240272 337878
rect 240232 334688 240284 334694
rect 240232 334630 240284 334636
rect 240336 330750 240364 338014
rect 240474 337770 240502 338028
rect 240566 337906 240594 338028
rect 240704 338014 240764 338042
rect 240566 337878 240640 337906
rect 240474 337742 240548 337770
rect 240324 330744 240376 330750
rect 240324 330686 240376 330692
rect 240048 326528 240100 326534
rect 240048 326470 240100 326476
rect 239404 326392 239456 326398
rect 239404 326334 239456 326340
rect 239312 4888 239364 4894
rect 239312 4830 239364 4836
rect 239220 3732 239272 3738
rect 239220 3674 239272 3680
rect 239324 480 239352 4830
rect 239416 3670 239444 326334
rect 240520 324970 240548 337742
rect 240612 333334 240640 337878
rect 240600 333328 240652 333334
rect 240600 333270 240652 333276
rect 240704 329254 240732 338014
rect 240842 337770 240870 338028
rect 240934 337906 240962 338028
rect 241072 338014 241132 338042
rect 240934 337878 241008 337906
rect 240842 337742 240916 337770
rect 240692 329248 240744 329254
rect 240692 329190 240744 329196
rect 240888 326602 240916 337742
rect 240980 333402 241008 337878
rect 240968 333396 241020 333402
rect 240968 333338 241020 333344
rect 241072 329322 241100 338014
rect 241210 337770 241238 338028
rect 241302 337906 241330 338028
rect 241440 338014 241500 338042
rect 241302 337878 241376 337906
rect 241164 337742 241238 337770
rect 241060 329316 241112 329322
rect 241060 329258 241112 329264
rect 240876 326596 240928 326602
rect 240876 326538 240928 326544
rect 240508 324964 240560 324970
rect 240508 324906 240560 324912
rect 241164 321554 241192 337742
rect 241348 332110 241376 337878
rect 241336 332104 241388 332110
rect 241336 332046 241388 332052
rect 241440 329390 241468 338014
rect 241578 337770 241606 338028
rect 241670 337906 241698 338028
rect 241808 338014 241868 338042
rect 241670 337878 241744 337906
rect 241578 337742 241652 337770
rect 241520 337680 241572 337686
rect 241520 337622 241572 337628
rect 241532 337278 241560 337622
rect 241520 337272 241572 337278
rect 241520 337214 241572 337220
rect 241428 329384 241480 329390
rect 241428 329326 241480 329332
rect 241624 326738 241652 337742
rect 241716 337210 241744 337878
rect 241704 337204 241756 337210
rect 241704 337146 241756 337152
rect 241808 330818 241836 338014
rect 241946 337770 241974 338028
rect 242038 337890 242066 338028
rect 242176 338014 242236 338042
rect 242026 337884 242078 337890
rect 242026 337826 242078 337832
rect 241946 337742 242112 337770
rect 241796 330812 241848 330818
rect 241796 330754 241848 330760
rect 241612 326732 241664 326738
rect 241612 326674 241664 326680
rect 242084 325038 242112 337742
rect 242176 329458 242204 338014
rect 242314 337770 242342 338028
rect 242268 337742 242342 337770
rect 242406 337770 242434 338028
rect 242498 337906 242526 338028
rect 242636 338014 242696 338042
rect 242498 337878 242572 337906
rect 242406 337742 242480 337770
rect 242164 329452 242216 329458
rect 242164 329394 242216 329400
rect 242268 325174 242296 337742
rect 242452 333470 242480 337742
rect 242440 333464 242492 333470
rect 242440 333406 242492 333412
rect 242544 329526 242572 337878
rect 242532 329520 242584 329526
rect 242532 329462 242584 329468
rect 242256 325168 242308 325174
rect 242256 325110 242308 325116
rect 242072 325032 242124 325038
rect 242072 324974 242124 324980
rect 242636 321554 242664 338014
rect 242774 337906 242802 338028
rect 242728 337878 242802 337906
rect 242728 331430 242756 337878
rect 242866 337770 242894 338028
rect 242820 337742 242894 337770
rect 243004 338014 243064 338042
rect 242716 331424 242768 331430
rect 242716 331366 242768 331372
rect 242820 330886 242848 337742
rect 242900 337680 242952 337686
rect 242900 337622 242952 337628
rect 242912 337346 242940 337622
rect 242900 337340 242952 337346
rect 242900 337282 242952 337288
rect 243004 334626 243032 338014
rect 243142 337770 243170 338028
rect 243234 337890 243262 338028
rect 243372 338014 243432 338042
rect 243372 337890 243400 338014
rect 243222 337884 243274 337890
rect 243222 337826 243274 337832
rect 243360 337884 243412 337890
rect 243360 337826 243412 337832
rect 243510 337770 243538 338028
rect 243602 337906 243630 338028
rect 243740 338014 243800 338042
rect 243602 337878 243676 337906
rect 243142 337742 243308 337770
rect 243084 337680 243136 337686
rect 243084 337622 243136 337628
rect 242992 334620 243044 334626
rect 242992 334562 243044 334568
rect 243096 331214 243124 337622
rect 243004 331186 243124 331214
rect 242808 330880 242860 330886
rect 242808 330822 242860 330828
rect 240520 321526 241192 321554
rect 241992 321526 242664 321554
rect 240520 11762 240548 321526
rect 240508 11756 240560 11762
rect 240508 11698 240560 11704
rect 240508 5432 240560 5438
rect 240508 5374 240560 5380
rect 239404 3664 239456 3670
rect 239404 3606 239456 3612
rect 240520 480 240548 5374
rect 241704 4684 241756 4690
rect 241704 4626 241756 4632
rect 241716 480 241744 4626
rect 241992 3942 242020 321526
rect 242900 4616 242952 4622
rect 242900 4558 242952 4564
rect 241980 3936 242032 3942
rect 241980 3878 242032 3884
rect 242912 480 242940 4558
rect 243004 4078 243032 331186
rect 243084 326460 243136 326466
rect 243084 326402 243136 326408
rect 242992 4072 243044 4078
rect 242992 4014 243044 4020
rect 243096 3398 243124 326402
rect 243176 326392 243228 326398
rect 243176 326334 243228 326340
rect 243188 4146 243216 326334
rect 243280 9042 243308 337742
rect 243372 337742 243538 337770
rect 243372 9110 243400 337742
rect 243648 334762 243676 337878
rect 243636 334756 243688 334762
rect 243636 334698 243688 334704
rect 243452 334620 243504 334626
rect 243452 334562 243504 334568
rect 243360 9104 243412 9110
rect 243360 9046 243412 9052
rect 243268 9036 243320 9042
rect 243268 8978 243320 8984
rect 243176 4140 243228 4146
rect 243176 4082 243228 4088
rect 243464 4010 243492 334562
rect 243740 326398 243768 338014
rect 243878 337770 243906 338028
rect 243970 337906 243998 338028
rect 244108 338014 244168 338042
rect 243970 337878 244044 337906
rect 243832 337742 243906 337770
rect 243832 337414 243860 337742
rect 243820 337408 243872 337414
rect 243820 337350 243872 337356
rect 244016 333606 244044 337878
rect 244004 333600 244056 333606
rect 244004 333542 244056 333548
rect 244108 326466 244136 338014
rect 244246 337770 244274 338028
rect 244338 337906 244366 338028
rect 244338 337878 244412 337906
rect 244200 337742 244274 337770
rect 244200 337482 244228 337742
rect 244188 337476 244240 337482
rect 244188 337418 244240 337424
rect 244384 329594 244412 337878
rect 244522 337770 244550 338028
rect 244614 337872 244642 338028
rect 244706 337940 244734 338028
rect 244844 338014 244904 338042
rect 244706 337912 244780 337940
rect 244614 337844 244688 337872
rect 244522 337742 244596 337770
rect 244372 329588 244424 329594
rect 244372 329530 244424 329536
rect 244096 326460 244148 326466
rect 244096 326402 244148 326408
rect 243728 326392 243780 326398
rect 243728 326334 243780 326340
rect 244096 4412 244148 4418
rect 244096 4354 244148 4360
rect 243452 4004 243504 4010
rect 243452 3946 243504 3952
rect 243084 3392 243136 3398
rect 243084 3334 243136 3340
rect 244108 480 244136 4354
rect 244568 3330 244596 337742
rect 244660 332178 244688 337844
rect 244648 332172 244700 332178
rect 244648 332114 244700 332120
rect 244752 327962 244780 337912
rect 244740 327956 244792 327962
rect 244740 327898 244792 327904
rect 244844 321554 244872 338014
rect 244982 337958 245010 338028
rect 244970 337952 245022 337958
rect 244970 337894 245022 337900
rect 245074 337822 245102 338028
rect 245212 338014 245272 338042
rect 245062 337816 245114 337822
rect 245062 337758 245114 337764
rect 245014 335472 245070 335481
rect 245014 335407 245070 335416
rect 244924 334620 244976 334626
rect 244924 334562 244976 334568
rect 244752 321526 244872 321554
rect 244556 3324 244608 3330
rect 244556 3266 244608 3272
rect 244752 3262 244780 321526
rect 244936 316034 244964 334562
rect 245028 331214 245056 335407
rect 245212 334626 245240 338014
rect 245350 337770 245378 338028
rect 245442 337906 245470 338028
rect 245580 338014 245640 338042
rect 245442 337878 245516 337906
rect 245304 337742 245378 337770
rect 245200 334620 245252 334626
rect 245200 334562 245252 334568
rect 245028 331186 245148 331214
rect 245120 328234 245148 331186
rect 245304 330954 245332 337742
rect 245488 336433 245516 337878
rect 245474 336424 245530 336433
rect 245474 336359 245530 336368
rect 245292 330948 245344 330954
rect 245292 330890 245344 330896
rect 245108 328228 245160 328234
rect 245108 328170 245160 328176
rect 245580 316034 245608 338014
rect 245718 337770 245746 338028
rect 245672 337742 245746 337770
rect 245810 337770 245838 338028
rect 245948 338014 246008 338042
rect 245810 337742 245884 337770
rect 245672 332246 245700 337742
rect 245752 337680 245804 337686
rect 245752 337622 245804 337628
rect 245660 332240 245712 332246
rect 245660 332182 245712 332188
rect 245764 331022 245792 337622
rect 245752 331016 245804 331022
rect 245752 330958 245804 330964
rect 245856 328030 245884 337742
rect 245844 328024 245896 328030
rect 245844 327966 245896 327972
rect 245948 325106 245976 338014
rect 246086 337958 246114 338028
rect 246074 337952 246126 337958
rect 246074 337894 246126 337900
rect 246178 337890 246206 338028
rect 246166 337884 246218 337890
rect 246166 337826 246218 337832
rect 246270 337770 246298 338028
rect 246224 337742 246298 337770
rect 246408 338014 246468 338042
rect 246028 337680 246080 337686
rect 246028 337622 246080 337628
rect 246040 328098 246068 337622
rect 246028 328092 246080 328098
rect 246028 328034 246080 328040
rect 246120 326392 246172 326398
rect 246120 326334 246172 326340
rect 245936 325100 245988 325106
rect 245936 325042 245988 325048
rect 244844 316006 244964 316034
rect 245120 316006 245608 316034
rect 244740 3256 244792 3262
rect 244740 3198 244792 3204
rect 244844 3194 244872 316006
rect 244832 3188 244884 3194
rect 244832 3130 244884 3136
rect 245120 3126 245148 316006
rect 245200 3460 245252 3466
rect 245200 3402 245252 3408
rect 245108 3120 245160 3126
rect 245108 3062 245160 3068
rect 245212 480 245240 3402
rect 246132 2990 246160 326334
rect 246224 3058 246252 337742
rect 246408 334626 246436 338014
rect 246546 337770 246574 338028
rect 246638 337958 246666 338028
rect 246776 338014 246836 338042
rect 246626 337952 246678 337958
rect 246626 337894 246678 337900
rect 246500 337742 246574 337770
rect 246396 334620 246448 334626
rect 246396 334562 246448 334568
rect 246500 331214 246528 337742
rect 246580 334620 246632 334626
rect 246580 334562 246632 334568
rect 246408 331186 246528 331214
rect 246408 328166 246436 331186
rect 246592 331090 246620 334562
rect 246580 331084 246632 331090
rect 246580 331026 246632 331032
rect 246396 328160 246448 328166
rect 246396 328102 246448 328108
rect 246776 316034 246804 338014
rect 246914 337770 246942 338028
rect 246868 337742 246942 337770
rect 246868 326670 246896 337742
rect 247006 337634 247034 338028
rect 247190 337770 247218 338028
rect 247282 337958 247310 338028
rect 247270 337952 247322 337958
rect 247270 337894 247322 337900
rect 247374 337906 247402 338028
rect 247512 338014 247572 338042
rect 247374 337878 247448 337906
rect 247316 337816 247368 337822
rect 247190 337742 247264 337770
rect 247316 337758 247368 337764
rect 246960 337606 247034 337634
rect 247132 337680 247184 337686
rect 247132 337622 247184 337628
rect 246856 326664 246908 326670
rect 246856 326606 246908 326612
rect 246960 326398 246988 337606
rect 247144 335481 247172 337622
rect 247130 335472 247186 335481
rect 247130 335407 247186 335416
rect 246948 326392 247000 326398
rect 246948 326334 247000 326340
rect 247132 326392 247184 326398
rect 247132 326334 247184 326340
rect 246408 316006 246804 316034
rect 246408 10334 246436 316006
rect 246396 10328 246448 10334
rect 246396 10270 246448 10276
rect 247144 5098 247172 326334
rect 247236 326262 247264 337742
rect 247224 326256 247276 326262
rect 247224 326198 247276 326204
rect 247224 326120 247276 326126
rect 247224 326062 247276 326068
rect 247236 6254 247264 326062
rect 247328 7682 247356 337758
rect 247420 326346 247448 337878
rect 247512 331214 247540 338014
rect 247650 337770 247678 338028
rect 247742 337958 247770 338028
rect 247880 338014 247940 338042
rect 247730 337952 247782 337958
rect 247730 337894 247782 337900
rect 247604 337742 247678 337770
rect 247604 332314 247632 337742
rect 247880 335889 247908 338014
rect 248018 337770 248046 338028
rect 248110 337822 248138 338028
rect 248248 338014 248308 338042
rect 247972 337742 248046 337770
rect 248098 337816 248150 337822
rect 248098 337758 248150 337764
rect 247866 335880 247922 335889
rect 247866 335815 247922 335824
rect 247972 334830 248000 337742
rect 247960 334824 248012 334830
rect 247960 334766 248012 334772
rect 247592 332308 247644 332314
rect 247592 332250 247644 332256
rect 247512 331186 247724 331214
rect 247420 326318 247632 326346
rect 247408 326256 247460 326262
rect 247408 326198 247460 326204
rect 247500 326256 247552 326262
rect 247500 326198 247552 326204
rect 247420 10402 247448 326198
rect 247512 10470 247540 326198
rect 247500 10464 247552 10470
rect 247500 10406 247552 10412
rect 247408 10396 247460 10402
rect 247408 10338 247460 10344
rect 247316 7676 247368 7682
rect 247316 7618 247368 7624
rect 247604 6914 247632 326318
rect 247696 326262 247724 331186
rect 248248 326398 248276 338014
rect 248386 337770 248414 338028
rect 248340 337742 248414 337770
rect 248478 337770 248506 338028
rect 248616 338014 248676 338042
rect 248478 337742 248552 337770
rect 248236 326392 248288 326398
rect 248236 326334 248288 326340
rect 247684 326256 247736 326262
rect 247684 326198 247736 326204
rect 248340 326126 248368 337742
rect 248524 328454 248552 337742
rect 248616 334898 248644 338014
rect 248754 337770 248782 338028
rect 248708 337742 248782 337770
rect 248846 337770 248874 338028
rect 248984 338014 249044 338042
rect 248846 337742 248920 337770
rect 248604 334892 248656 334898
rect 248604 334834 248656 334840
rect 248708 333674 248736 337742
rect 248696 333668 248748 333674
rect 248696 333610 248748 333616
rect 248892 328454 248920 337742
rect 248984 334966 249012 338014
rect 249122 337906 249150 338028
rect 249076 337878 249150 337906
rect 248972 334960 249024 334966
rect 248972 334902 249024 334908
rect 249076 332382 249104 337878
rect 249214 337770 249242 338028
rect 249168 337742 249242 337770
rect 249352 338014 249412 338042
rect 249064 332376 249116 332382
rect 249064 332318 249116 332324
rect 248524 328426 248828 328454
rect 248892 328426 249012 328454
rect 248696 326392 248748 326398
rect 248696 326334 248748 326340
rect 248328 326120 248380 326126
rect 248328 326062 248380 326068
rect 248708 9246 248736 326334
rect 248696 9240 248748 9246
rect 248696 9182 248748 9188
rect 248800 7750 248828 328426
rect 248984 9178 249012 328426
rect 249168 326398 249196 337742
rect 249352 335102 249380 338014
rect 249490 337770 249518 338028
rect 249444 337742 249518 337770
rect 249582 337770 249610 338028
rect 249720 338014 249780 338042
rect 249582 337742 249656 337770
rect 249340 335096 249392 335102
rect 249340 335038 249392 335044
rect 249444 332450 249472 337742
rect 249432 332444 249484 332450
rect 249432 332386 249484 332392
rect 249156 326392 249208 326398
rect 249156 326334 249208 326340
rect 249628 316034 249656 337742
rect 249720 335170 249748 338014
rect 249858 337770 249886 338028
rect 249812 337742 249886 337770
rect 249950 337770 249978 338028
rect 250042 337906 250070 338028
rect 250180 338014 250240 338042
rect 250042 337878 250116 337906
rect 249950 337742 250024 337770
rect 249708 335164 249760 335170
rect 249708 335106 249760 335112
rect 249812 333742 249840 337742
rect 249800 333736 249852 333742
rect 249800 333678 249852 333684
rect 249996 329730 250024 337742
rect 250088 335238 250116 337878
rect 250076 335232 250128 335238
rect 250076 335174 250128 335180
rect 250180 332518 250208 338014
rect 250318 337770 250346 338028
rect 250410 337872 250438 338028
rect 250548 338014 250608 338042
rect 250410 337844 250484 337872
rect 250272 337742 250346 337770
rect 250168 332512 250220 332518
rect 250168 332454 250220 332460
rect 249984 329724 250036 329730
rect 249984 329666 250036 329672
rect 250272 316034 250300 337742
rect 250456 335306 250484 337844
rect 250444 335300 250496 335306
rect 250444 335242 250496 335248
rect 250548 332586 250576 338014
rect 250686 337770 250714 338028
rect 250778 337906 250806 338028
rect 250916 338014 250976 338042
rect 250778 337878 250852 337906
rect 250640 337742 250714 337770
rect 250536 332580 250588 332586
rect 250536 332522 250588 332528
rect 250640 331158 250668 337742
rect 250720 337680 250772 337686
rect 250720 337622 250772 337628
rect 250732 331838 250760 337622
rect 250824 334558 250852 337878
rect 250916 337822 250944 338014
rect 250904 337816 250956 337822
rect 250904 337758 250956 337764
rect 250904 337680 250956 337686
rect 251054 337634 251082 338028
rect 251146 337958 251174 338028
rect 251284 338014 251344 338042
rect 251134 337952 251186 337958
rect 251134 337894 251186 337900
rect 250904 337622 250956 337628
rect 250812 334552 250864 334558
rect 250812 334494 250864 334500
rect 250916 334490 250944 337622
rect 251008 337606 251082 337634
rect 250904 334484 250956 334490
rect 250904 334426 250956 334432
rect 250720 331832 250772 331838
rect 250720 331774 250772 331780
rect 250628 331152 250680 331158
rect 250628 331094 250680 331100
rect 251008 316034 251036 337606
rect 251284 336190 251312 338014
rect 251422 337770 251450 338028
rect 251514 337890 251542 338028
rect 251502 337884 251554 337890
rect 251502 337826 251554 337832
rect 251698 337770 251726 338028
rect 251790 337890 251818 338028
rect 251882 337906 251910 338028
rect 252020 338014 252080 338042
rect 251778 337884 251830 337890
rect 251882 337878 251956 337906
rect 251778 337826 251830 337832
rect 251422 337742 251496 337770
rect 251698 337742 251864 337770
rect 251468 336274 251496 337742
rect 251732 337680 251784 337686
rect 251732 337622 251784 337628
rect 251468 336246 251588 336274
rect 251272 336184 251324 336190
rect 251272 336126 251324 336132
rect 251456 336184 251508 336190
rect 251456 336126 251508 336132
rect 251364 323060 251416 323066
rect 251364 323002 251416 323008
rect 249260 316006 249656 316034
rect 250180 316006 250300 316034
rect 250364 316006 251036 316034
rect 249260 9314 249288 316006
rect 250180 10538 250208 316006
rect 250364 17270 250392 316006
rect 250352 17264 250404 17270
rect 250352 17206 250404 17212
rect 250168 10532 250220 10538
rect 250168 10474 250220 10480
rect 249248 9308 249300 9314
rect 249248 9250 249300 9256
rect 248972 9172 249024 9178
rect 248972 9114 249024 9120
rect 251376 7886 251404 323002
rect 251364 7880 251416 7886
rect 251364 7822 251416 7828
rect 251468 7818 251496 336126
rect 251560 9382 251588 336246
rect 251640 334620 251692 334626
rect 251640 334562 251692 334568
rect 251548 9376 251600 9382
rect 251548 9318 251600 9324
rect 251652 8022 251680 334562
rect 251744 323066 251772 337622
rect 251836 336274 251864 337742
rect 251928 336734 251956 337878
rect 251916 336728 251968 336734
rect 251916 336670 251968 336676
rect 251836 336246 251956 336274
rect 251824 336184 251876 336190
rect 251824 336126 251876 336132
rect 251732 323060 251784 323066
rect 251732 323002 251784 323008
rect 251640 8016 251692 8022
rect 251640 7958 251692 7964
rect 251456 7812 251508 7818
rect 251456 7754 251508 7760
rect 248788 7744 248840 7750
rect 248788 7686 248840 7692
rect 247512 6886 247632 6914
rect 247224 6248 247276 6254
rect 247224 6190 247276 6196
rect 247132 5092 247184 5098
rect 247132 5034 247184 5040
rect 246396 4480 246448 4486
rect 246396 4422 246448 4428
rect 246212 3052 246264 3058
rect 246212 2994 246264 3000
rect 246120 2984 246172 2990
rect 246120 2926 246172 2932
rect 246408 480 246436 4422
rect 247512 2922 247540 6886
rect 249984 4752 250036 4758
rect 249984 4694 250036 4700
rect 247592 4548 247644 4554
rect 247592 4490 247644 4496
rect 247500 2916 247552 2922
rect 247500 2858 247552 2864
rect 247604 480 247632 4490
rect 248788 3936 248840 3942
rect 248788 3878 248840 3884
rect 248800 480 248828 3878
rect 249996 480 250024 4694
rect 251836 4418 251864 336126
rect 251928 333810 251956 336246
rect 252020 333878 252048 338014
rect 252158 337770 252186 338028
rect 252112 337742 252186 337770
rect 252250 337770 252278 338028
rect 252388 338014 252448 338042
rect 252250 337742 252324 337770
rect 252008 333872 252060 333878
rect 252008 333814 252060 333820
rect 251916 333804 251968 333810
rect 251916 333746 251968 333752
rect 252112 316034 252140 337742
rect 252296 335578 252324 337742
rect 252284 335572 252336 335578
rect 252284 335514 252336 335520
rect 252388 333198 252416 338014
rect 252526 337770 252554 338028
rect 252480 337742 252554 337770
rect 252480 334626 252508 337742
rect 252618 337736 252646 338028
rect 252756 338014 252816 338042
rect 252618 337708 252692 337736
rect 252664 337634 252692 337708
rect 252572 337606 252692 337634
rect 252572 336462 252600 337606
rect 252560 336456 252612 336462
rect 252560 336398 252612 336404
rect 252652 336456 252704 336462
rect 252652 336398 252704 336404
rect 252560 336252 252612 336258
rect 252560 336194 252612 336200
rect 252468 334620 252520 334626
rect 252468 334562 252520 334568
rect 252572 334422 252600 336194
rect 252560 334416 252612 334422
rect 252560 334358 252612 334364
rect 252376 333192 252428 333198
rect 252376 333134 252428 333140
rect 252664 332926 252692 336398
rect 252652 332920 252704 332926
rect 252652 332862 252704 332868
rect 252020 316006 252140 316034
rect 252020 7954 252048 316006
rect 252008 7948 252060 7954
rect 252008 7890 252060 7896
rect 252756 6322 252784 338014
rect 252894 337770 252922 338028
rect 252986 337906 253014 338028
rect 253124 338014 253184 338042
rect 252986 337878 253060 337906
rect 253124 337890 253152 338014
rect 253262 337906 253290 338028
rect 252894 337742 252968 337770
rect 252836 334620 252888 334626
rect 252836 334562 252888 334568
rect 252848 6526 252876 334562
rect 252940 325106 252968 337742
rect 253032 336054 253060 337878
rect 253112 337884 253164 337890
rect 253112 337826 253164 337832
rect 253216 337878 253290 337906
rect 253112 337748 253164 337754
rect 253112 337690 253164 337696
rect 253020 336048 253072 336054
rect 253020 335990 253072 335996
rect 252928 325100 252980 325106
rect 252928 325042 252980 325048
rect 253020 324896 253072 324902
rect 253020 324838 253072 324844
rect 252928 319320 252980 319326
rect 252928 319262 252980 319268
rect 252940 8158 252968 319262
rect 252928 8152 252980 8158
rect 252928 8094 252980 8100
rect 253032 8090 253060 324838
rect 253124 319326 253152 337690
rect 253112 319320 253164 319326
rect 253112 319262 253164 319268
rect 253216 316034 253244 337878
rect 253354 337770 253382 338028
rect 253308 337742 253382 337770
rect 253538 337770 253566 338028
rect 253630 337890 253658 338028
rect 253722 337890 253750 338028
rect 253618 337884 253670 337890
rect 253618 337826 253670 337832
rect 253710 337884 253762 337890
rect 253710 337826 253762 337832
rect 253814 337770 253842 338028
rect 253538 337742 253704 337770
rect 253308 335442 253336 337742
rect 253388 337680 253440 337686
rect 253388 337622 253440 337628
rect 253572 337680 253624 337686
rect 253572 337622 253624 337628
rect 253296 335436 253348 335442
rect 253296 335378 253348 335384
rect 253124 316006 253244 316034
rect 253020 8084 253072 8090
rect 253020 8026 253072 8032
rect 253124 7614 253152 316006
rect 253112 7608 253164 7614
rect 253112 7550 253164 7556
rect 252836 6520 252888 6526
rect 252836 6462 252888 6468
rect 253400 6458 253428 337622
rect 253584 336734 253612 337622
rect 253572 336728 253624 336734
rect 253572 336670 253624 336676
rect 253388 6452 253440 6458
rect 253388 6394 253440 6400
rect 253676 6390 253704 337742
rect 253768 337742 253842 337770
rect 253952 338014 254012 338042
rect 253768 334626 253796 337742
rect 253848 335572 253900 335578
rect 253848 335514 253900 335520
rect 253756 334620 253808 334626
rect 253756 334562 253808 334568
rect 253664 6384 253716 6390
rect 253664 6326 253716 6332
rect 252744 6316 252796 6322
rect 252744 6258 252796 6264
rect 253860 5506 253888 335514
rect 253952 331770 253980 338014
rect 254090 337770 254118 338028
rect 254182 337906 254210 338028
rect 254320 338014 254380 338042
rect 254182 337878 254256 337906
rect 254044 337742 254118 337770
rect 254044 336122 254072 337742
rect 254032 336116 254084 336122
rect 254032 336058 254084 336064
rect 254228 333946 254256 337878
rect 254216 333940 254268 333946
rect 254216 333882 254268 333888
rect 253940 331764 253992 331770
rect 253940 331706 253992 331712
rect 254320 331702 254348 338014
rect 254458 337770 254486 338028
rect 254550 337906 254578 338028
rect 254688 338014 254748 338042
rect 254550 337878 254624 337906
rect 254412 337742 254486 337770
rect 254412 335646 254440 337742
rect 254400 335640 254452 335646
rect 254400 335582 254452 335588
rect 254596 333130 254624 337878
rect 254584 333124 254636 333130
rect 254584 333066 254636 333072
rect 254584 332988 254636 332994
rect 254584 332930 254636 332936
rect 254308 331696 254360 331702
rect 254308 331638 254360 331644
rect 253480 5500 253532 5506
rect 253480 5442 253532 5448
rect 253848 5500 253900 5506
rect 253848 5442 253900 5448
rect 251824 4412 251876 4418
rect 251824 4354 251876 4360
rect 251180 4072 251232 4078
rect 251180 4014 251232 4020
rect 251192 480 251220 4014
rect 252376 3596 252428 3602
rect 252376 3538 252428 3544
rect 252388 480 252416 3538
rect 253492 480 253520 5442
rect 254596 5030 254624 332930
rect 254688 331226 254716 338014
rect 254826 337770 254854 338028
rect 254780 337742 254854 337770
rect 254780 335918 254808 337742
rect 254918 337668 254946 338028
rect 254872 337640 254946 337668
rect 255056 338014 255116 338042
rect 254768 335912 254820 335918
rect 254768 335854 254820 335860
rect 254872 335764 254900 337640
rect 254780 335736 254900 335764
rect 254780 334286 254808 335736
rect 254860 335368 254912 335374
rect 254860 335310 254912 335316
rect 254768 334280 254820 334286
rect 254768 334222 254820 334228
rect 254676 331220 254728 331226
rect 254676 331162 254728 331168
rect 254872 330410 254900 335310
rect 255056 330478 255084 338014
rect 255194 337770 255222 338028
rect 255148 337742 255222 337770
rect 255148 335850 255176 337742
rect 255286 337668 255314 338028
rect 255240 337640 255314 337668
rect 255424 338014 255484 338042
rect 255136 335844 255188 335850
rect 255136 335786 255188 335792
rect 255240 333062 255268 337640
rect 255228 333056 255280 333062
rect 255228 332998 255280 333004
rect 255424 330478 255452 338014
rect 255562 337770 255590 338028
rect 255654 337822 255682 338028
rect 255792 338014 255852 338042
rect 255516 337742 255590 337770
rect 255642 337816 255694 337822
rect 255642 337758 255694 337764
rect 255044 330472 255096 330478
rect 255044 330414 255096 330420
rect 255412 330472 255464 330478
rect 255412 330414 255464 330420
rect 254860 330404 254912 330410
rect 254860 330346 254912 330352
rect 255412 330268 255464 330274
rect 255412 330210 255464 330216
rect 255424 5370 255452 330210
rect 255412 5364 255464 5370
rect 255412 5306 255464 5312
rect 255516 5166 255544 337742
rect 255688 337680 255740 337686
rect 255688 337622 255740 337628
rect 255596 330540 255648 330546
rect 255596 330482 255648 330488
rect 255608 5302 255636 330482
rect 255700 6662 255728 337622
rect 255792 335374 255820 338014
rect 255930 337770 255958 338028
rect 256022 337890 256050 338028
rect 256160 338014 256220 338042
rect 256010 337884 256062 337890
rect 256010 337826 256062 337832
rect 255930 337742 256004 337770
rect 255780 335368 255832 335374
rect 255780 335310 255832 335316
rect 255976 330562 256004 337742
rect 256160 336462 256188 338014
rect 256298 337770 256326 338028
rect 256252 337742 256326 337770
rect 256148 336456 256200 336462
rect 256148 336398 256200 336404
rect 255976 330534 256096 330562
rect 256252 330546 256280 337742
rect 256390 337668 256418 338028
rect 256344 337640 256418 337668
rect 256528 338014 256588 338042
rect 255964 330472 256016 330478
rect 255964 330414 256016 330420
rect 255780 330336 255832 330342
rect 255780 330278 255832 330284
rect 255872 330336 255924 330342
rect 255872 330278 255924 330284
rect 255688 6656 255740 6662
rect 255688 6598 255740 6604
rect 255792 6594 255820 330278
rect 255884 6730 255912 330278
rect 255976 8226 256004 330414
rect 255964 8220 256016 8226
rect 255964 8162 256016 8168
rect 255872 6724 255924 6730
rect 255872 6666 255924 6672
rect 255780 6588 255832 6594
rect 255780 6530 255832 6536
rect 255596 5296 255648 5302
rect 255596 5238 255648 5244
rect 256068 5234 256096 330534
rect 256240 330540 256292 330546
rect 256240 330482 256292 330488
rect 256344 330342 256372 337640
rect 256528 332858 256556 338014
rect 256666 337770 256694 338028
rect 256758 337906 256786 338028
rect 256896 338014 256956 338042
rect 256758 337878 256832 337906
rect 256620 337742 256694 337770
rect 256516 332852 256568 332858
rect 256516 332794 256568 332800
rect 256332 330336 256384 330342
rect 256332 330278 256384 330284
rect 256620 330274 256648 337742
rect 256804 334218 256832 337878
rect 256792 334212 256844 334218
rect 256792 334154 256844 334160
rect 256896 331634 256924 338014
rect 257034 337770 257062 338028
rect 257126 337906 257154 338028
rect 257264 338014 257324 338042
rect 257126 337878 257200 337906
rect 256988 337742 257062 337770
rect 256988 336394 257016 337742
rect 256976 336388 257028 336394
rect 256976 336330 257028 336336
rect 257172 332790 257200 337878
rect 257160 332784 257212 332790
rect 257160 332726 257212 332732
rect 256884 331628 256936 331634
rect 256884 331570 256936 331576
rect 257264 330410 257292 338014
rect 257402 337770 257430 338028
rect 257356 337742 257430 337770
rect 257494 337770 257522 338028
rect 257586 337906 257614 338028
rect 257724 338014 257784 338042
rect 257586 337878 257660 337906
rect 257494 337742 257568 337770
rect 257356 335510 257384 337742
rect 257436 337680 257488 337686
rect 257436 337622 257488 337628
rect 257344 335504 257396 335510
rect 257344 335446 257396 335452
rect 257344 334756 257396 334762
rect 257344 334698 257396 334704
rect 257252 330404 257304 330410
rect 257252 330346 257304 330352
rect 256608 330268 256660 330274
rect 256608 330210 256660 330216
rect 256056 5228 256108 5234
rect 256056 5170 256108 5176
rect 255504 5160 255556 5166
rect 255504 5102 255556 5108
rect 254584 5024 254636 5030
rect 254584 4966 254636 4972
rect 257068 4140 257120 4146
rect 257068 4082 257120 4088
rect 255872 3800 255924 3806
rect 255872 3742 255924 3748
rect 254676 3732 254728 3738
rect 254676 3674 254728 3680
rect 254688 480 254716 3674
rect 255884 480 255912 3742
rect 257080 480 257108 4082
rect 257356 3466 257384 334698
rect 257448 9450 257476 337622
rect 257540 334150 257568 337742
rect 257528 334144 257580 334150
rect 257528 334086 257580 334092
rect 257632 330206 257660 337878
rect 257724 335442 257752 338014
rect 257862 337770 257890 338028
rect 257954 337906 257982 338028
rect 258092 338014 258152 338042
rect 257954 337878 258028 337906
rect 257816 337742 257890 337770
rect 257712 335436 257764 335442
rect 257712 335378 257764 335384
rect 257816 332722 257844 337742
rect 257804 332716 257856 332722
rect 257804 332658 257856 332664
rect 258000 331566 258028 337878
rect 258092 336530 258120 338014
rect 258230 337770 258258 338028
rect 258184 337742 258258 337770
rect 258080 336524 258132 336530
rect 258080 336466 258132 336472
rect 258184 332654 258212 337742
rect 258322 337736 258350 338028
rect 258460 338014 258520 338042
rect 258322 337708 258396 337736
rect 258368 337668 258396 337708
rect 258276 337640 258396 337668
rect 258276 334082 258304 337640
rect 258460 335782 258488 338014
rect 258598 337770 258626 338028
rect 258690 337822 258718 338028
rect 258828 338014 258888 338042
rect 258552 337742 258626 337770
rect 258678 337816 258730 337822
rect 258678 337758 258730 337764
rect 258448 335776 258500 335782
rect 258448 335718 258500 335724
rect 258356 334620 258408 334626
rect 258356 334562 258408 334568
rect 258264 334076 258316 334082
rect 258264 334018 258316 334024
rect 258172 332648 258224 332654
rect 258172 332590 258224 332596
rect 257988 331560 258040 331566
rect 257988 331502 258040 331508
rect 257620 330200 257672 330206
rect 257620 330142 257672 330148
rect 257436 9444 257488 9450
rect 257436 9386 257488 9392
rect 258368 4962 258396 334562
rect 258552 334014 258580 337742
rect 258828 336258 258856 338014
rect 258966 337770 258994 338028
rect 259058 337906 259086 338028
rect 259196 338014 259256 338042
rect 259058 337878 259132 337906
rect 258920 337742 258994 337770
rect 258816 336252 258868 336258
rect 258816 336194 258868 336200
rect 258724 335368 258776 335374
rect 258724 335310 258776 335316
rect 258540 334008 258592 334014
rect 258540 333950 258592 333956
rect 258632 330540 258684 330546
rect 258632 330482 258684 330488
rect 258356 4956 258408 4962
rect 258356 4898 258408 4904
rect 258644 4826 258672 330482
rect 258736 5438 258764 335310
rect 258816 333260 258868 333266
rect 258816 333202 258868 333208
rect 258724 5432 258776 5438
rect 258724 5374 258776 5380
rect 258632 4820 258684 4826
rect 258632 4762 258684 4768
rect 258828 4690 258856 333202
rect 258920 331498 258948 337742
rect 259104 332994 259132 337878
rect 259196 335714 259224 338014
rect 259334 337770 259362 338028
rect 259288 337742 259362 337770
rect 259184 335708 259236 335714
rect 259184 335650 259236 335656
rect 259092 332988 259144 332994
rect 259092 332930 259144 332936
rect 258908 331492 258960 331498
rect 258908 331434 258960 331440
rect 259288 330546 259316 337742
rect 259426 337668 259454 338028
rect 259610 337770 259638 338028
rect 259702 337872 259730 338028
rect 259794 337940 259822 338028
rect 259932 338014 259992 338042
rect 259794 337912 259868 337940
rect 259702 337844 259776 337872
rect 259610 337742 259684 337770
rect 259380 337640 259454 337668
rect 259380 334626 259408 337640
rect 259368 334620 259420 334626
rect 259368 334562 259420 334568
rect 259656 330562 259684 337742
rect 259748 335374 259776 337844
rect 259736 335368 259788 335374
rect 259736 335310 259788 335316
rect 259840 333266 259868 337912
rect 259828 333260 259880 333266
rect 259828 333202 259880 333208
rect 259932 330562 259960 338014
rect 260070 337770 260098 338028
rect 260024 337742 260098 337770
rect 260024 336190 260052 337742
rect 260162 337668 260190 338028
rect 260116 337640 260190 337668
rect 260300 338014 260360 338042
rect 260012 336184 260064 336190
rect 260012 336126 260064 336132
rect 260116 336036 260144 337640
rect 260024 336008 260144 336036
rect 260024 334762 260052 336008
rect 260104 335504 260156 335510
rect 260104 335446 260156 335452
rect 260012 334756 260064 334762
rect 260012 334698 260064 334704
rect 260012 334620 260064 334626
rect 260012 334562 260064 334568
rect 259276 330540 259328 330546
rect 259656 330534 259776 330562
rect 259276 330482 259328 330488
rect 259644 330472 259696 330478
rect 259644 330414 259696 330420
rect 258816 4684 258868 4690
rect 258816 4626 258868 4632
rect 259656 4486 259684 330414
rect 259748 4894 259776 330534
rect 259840 330534 259960 330562
rect 259736 4888 259788 4894
rect 259736 4830 259788 4836
rect 259840 4622 259868 330534
rect 260024 316034 260052 334562
rect 259932 316006 260052 316034
rect 259828 4616 259880 4622
rect 259828 4558 259880 4564
rect 259644 4480 259696 4486
rect 259644 4422 259696 4428
rect 259932 4078 259960 316006
rect 260116 4146 260144 335446
rect 260300 330478 260328 338014
rect 260438 337872 260466 338028
rect 260392 337844 260466 337872
rect 260392 335986 260420 337844
rect 260530 337770 260558 338028
rect 260484 337742 260558 337770
rect 260668 338014 260728 338042
rect 260380 335980 260432 335986
rect 260380 335922 260432 335928
rect 260288 330472 260340 330478
rect 260288 330414 260340 330420
rect 260484 316034 260512 337742
rect 260668 336666 260696 338014
rect 260806 337906 260834 338028
rect 260760 337878 260834 337906
rect 260898 337906 260926 338028
rect 261036 338014 261096 338042
rect 260898 337878 260972 337906
rect 260656 336660 260708 336666
rect 260656 336602 260708 336608
rect 260656 335436 260708 335442
rect 260656 335378 260708 335384
rect 260668 331214 260696 335378
rect 260760 334626 260788 337878
rect 260840 337816 260892 337822
rect 260840 337758 260892 337764
rect 260748 334620 260800 334626
rect 260748 334562 260800 334568
rect 260668 331186 260788 331214
rect 260208 316006 260512 316034
rect 260104 4140 260156 4146
rect 260104 4082 260156 4088
rect 259920 4072 259972 4078
rect 259920 4014 259972 4020
rect 260208 3942 260236 316006
rect 260760 6914 260788 331186
rect 260852 330426 260880 337758
rect 260944 336444 260972 337878
rect 261036 336598 261064 338014
rect 261174 337770 261202 338028
rect 261266 337890 261294 338028
rect 261254 337884 261306 337890
rect 261254 337826 261306 337832
rect 261358 337770 261386 338028
rect 261174 337742 261248 337770
rect 261024 336592 261076 336598
rect 261024 336534 261076 336540
rect 260944 336416 261064 336444
rect 260852 330398 260972 330426
rect 260840 330336 260892 330342
rect 260840 330278 260892 330284
rect 260668 6886 260788 6914
rect 260196 3936 260248 3942
rect 260196 3878 260248 3884
rect 259460 3528 259512 3534
rect 259460 3470 259512 3476
rect 257344 3460 257396 3466
rect 257344 3402 257396 3408
rect 258264 3188 258316 3194
rect 258264 3130 258316 3136
rect 258276 480 258304 3130
rect 259472 480 259500 3470
rect 260668 480 260696 6886
rect 260852 3074 260880 330278
rect 260944 3806 260972 330398
rect 260932 3800 260984 3806
rect 260932 3742 260984 3748
rect 261036 3602 261064 336416
rect 261116 335368 261168 335374
rect 261116 335310 261168 335316
rect 261128 330342 261156 335310
rect 261116 330336 261168 330342
rect 261116 330278 261168 330284
rect 261116 330200 261168 330206
rect 261116 330142 261168 330148
rect 261024 3596 261076 3602
rect 261024 3538 261076 3544
rect 261128 3534 261156 330142
rect 261220 3738 261248 337742
rect 261312 337742 261386 337770
rect 261496 338014 261556 338042
rect 261312 335510 261340 337742
rect 261300 335504 261352 335510
rect 261300 335446 261352 335452
rect 261496 316034 261524 338014
rect 261634 337770 261662 338028
rect 261726 337906 261754 338028
rect 261864 338014 261924 338042
rect 261726 337878 261800 337906
rect 261588 337742 261662 337770
rect 261588 330206 261616 337742
rect 261772 335442 261800 337878
rect 261760 335436 261812 335442
rect 261760 335378 261812 335384
rect 261864 335374 261892 338014
rect 262002 337770 262030 338028
rect 262094 337906 262122 338028
rect 262232 338014 262292 338042
rect 262094 337878 262168 337906
rect 262002 337742 262076 337770
rect 261852 335368 261904 335374
rect 261852 335310 261904 335316
rect 261576 330200 261628 330206
rect 261576 330142 261628 330148
rect 262048 325694 262076 337742
rect 262140 335238 262168 337878
rect 262232 336462 262260 338014
rect 262370 337770 262398 338028
rect 262462 337872 262490 338028
rect 262600 338014 262660 338042
rect 262462 337844 262536 337872
rect 262370 337742 262444 337770
rect 262312 336660 262364 336666
rect 262312 336602 262364 336608
rect 262220 336456 262272 336462
rect 262220 336398 262272 336404
rect 262324 335578 262352 336602
rect 262312 335572 262364 335578
rect 262312 335514 262364 335520
rect 262128 335232 262180 335238
rect 262128 335174 262180 335180
rect 262416 334422 262444 337742
rect 262508 336666 262536 337844
rect 262496 336660 262548 336666
rect 262496 336602 262548 336608
rect 262496 336524 262548 336530
rect 262496 336466 262548 336472
rect 262404 334416 262456 334422
rect 262404 334358 262456 334364
rect 262048 325666 262168 325694
rect 261312 316006 261524 316034
rect 261208 3732 261260 3738
rect 261208 3674 261260 3680
rect 261116 3528 261168 3534
rect 261116 3470 261168 3476
rect 261312 3194 261340 316006
rect 262140 3534 262168 325666
rect 262508 5370 262536 336466
rect 262600 335442 262628 338014
rect 262738 337770 262766 338028
rect 262830 337872 262858 338028
rect 262968 338014 263028 338042
rect 262968 337958 262996 338014
rect 262956 337952 263008 337958
rect 262956 337894 263008 337900
rect 262830 337844 262904 337872
rect 262738 337742 262812 337770
rect 262784 335510 262812 337742
rect 262876 335730 262904 337844
rect 263106 337770 263134 338028
rect 263198 337906 263226 338028
rect 263336 338014 263396 338042
rect 263198 337878 263272 337906
rect 262968 337742 263134 337770
rect 262968 335918 262996 337742
rect 263048 337680 263100 337686
rect 263048 337622 263100 337628
rect 263060 336122 263088 337622
rect 263048 336116 263100 336122
rect 263048 336058 263100 336064
rect 262956 335912 263008 335918
rect 262956 335854 263008 335860
rect 262876 335702 262996 335730
rect 262772 335504 262824 335510
rect 262772 335446 262824 335452
rect 262588 335436 262640 335442
rect 262588 335378 262640 335384
rect 262864 335232 262916 335238
rect 262864 335174 262916 335180
rect 262496 5364 262548 5370
rect 262496 5306 262548 5312
rect 262128 3528 262180 3534
rect 262128 3470 262180 3476
rect 262876 3466 262904 335174
rect 262968 4690 262996 335702
rect 263244 334778 263272 337878
rect 263060 334750 263272 334778
rect 263060 4758 263088 334750
rect 263336 334642 263364 338014
rect 263474 337872 263502 338028
rect 263428 337844 263502 337872
rect 263428 336734 263456 337844
rect 263566 337770 263594 338028
rect 263520 337742 263594 337770
rect 263750 337770 263778 338028
rect 263842 337958 263870 338028
rect 263830 337952 263882 337958
rect 263934 337940 263962 338028
rect 263934 337912 264008 337940
rect 263830 337894 263882 337900
rect 263750 337742 263824 337770
rect 263520 336818 263548 337742
rect 263520 336790 263640 336818
rect 263416 336728 263468 336734
rect 263416 336670 263468 336676
rect 263612 336530 263640 336790
rect 263600 336524 263652 336530
rect 263600 336466 263652 336472
rect 263508 335504 263560 335510
rect 263508 335446 263560 335452
rect 263416 335436 263468 335442
rect 263416 335378 263468 335384
rect 263152 334614 263364 334642
rect 263152 5438 263180 334614
rect 263428 334506 263456 335378
rect 263244 334478 263456 334506
rect 263244 325694 263272 334478
rect 263416 334416 263468 334422
rect 263416 334358 263468 334364
rect 263244 325666 263364 325694
rect 263140 5432 263192 5438
rect 263140 5374 263192 5380
rect 263048 4752 263100 4758
rect 263048 4694 263100 4700
rect 262956 4684 263008 4690
rect 262956 4626 263008 4632
rect 262956 3528 263008 3534
rect 262956 3470 263008 3476
rect 262864 3460 262916 3466
rect 262864 3402 262916 3408
rect 261300 3188 261352 3194
rect 261300 3130 261352 3136
rect 260852 3046 261800 3074
rect 261772 480 261800 3046
rect 262968 480 262996 3470
rect 263336 3058 263364 325666
rect 263428 3602 263456 334358
rect 263416 3596 263468 3602
rect 263416 3538 263468 3544
rect 263520 3194 263548 335446
rect 263796 334422 263824 337742
rect 263876 336456 263928 336462
rect 263876 336398 263928 336404
rect 263784 334416 263836 334422
rect 263784 334358 263836 334364
rect 263888 330206 263916 336398
rect 263980 335730 264008 337912
rect 264118 337770 264146 338028
rect 264210 337958 264238 338028
rect 264198 337952 264250 337958
rect 264302 337940 264330 338028
rect 264440 338014 264500 338042
rect 264302 337912 264376 337940
rect 264198 337894 264250 337900
rect 264118 337742 264192 337770
rect 263980 335702 264100 335730
rect 263968 335028 264020 335034
rect 263968 334970 264020 334976
rect 263876 330200 263928 330206
rect 263876 330142 263928 330148
rect 263980 325694 264008 334970
rect 264072 333266 264100 335702
rect 264060 333260 264112 333266
rect 264060 333202 264112 333208
rect 264164 330290 264192 337742
rect 264348 334642 264376 337912
rect 264440 334778 264468 338014
rect 264578 337958 264606 338028
rect 264566 337952 264618 337958
rect 264670 337940 264698 338028
rect 264808 338014 264868 338042
rect 264670 337912 264744 337940
rect 264566 337894 264618 337900
rect 264716 337770 264744 337912
rect 264808 337890 264836 338014
rect 264796 337884 264848 337890
rect 264796 337826 264848 337832
rect 264946 337770 264974 338028
rect 264716 337742 264836 337770
rect 264704 337680 264756 337686
rect 264704 337622 264756 337628
rect 264716 336734 264744 337622
rect 264704 336728 264756 336734
rect 264704 336670 264756 336676
rect 264808 335034 264836 337742
rect 264900 337742 264974 337770
rect 265038 337770 265066 338028
rect 265130 337906 265158 338028
rect 265268 338014 265328 338042
rect 265130 337878 265204 337906
rect 265038 337742 265112 337770
rect 264796 335028 264848 335034
rect 264796 334970 264848 334976
rect 264440 334750 264744 334778
rect 264348 334614 264652 334642
rect 264244 334416 264296 334422
rect 264244 334358 264296 334364
rect 264256 330426 264284 334358
rect 264520 333260 264572 333266
rect 264520 333202 264572 333208
rect 264256 330398 264468 330426
rect 264164 330262 264376 330290
rect 264244 330200 264296 330206
rect 264244 330142 264296 330148
rect 263980 325666 264192 325694
rect 264164 4894 264192 325666
rect 264152 4888 264204 4894
rect 264152 4830 264204 4836
rect 264256 3534 264284 330142
rect 264348 5166 264376 330262
rect 264440 5302 264468 330398
rect 264428 5296 264480 5302
rect 264428 5238 264480 5244
rect 264532 5234 264560 333202
rect 264520 5228 264572 5234
rect 264520 5170 264572 5176
rect 264336 5160 264388 5166
rect 264336 5102 264388 5108
rect 264624 5098 264652 334614
rect 264612 5092 264664 5098
rect 264612 5034 264664 5040
rect 264716 5030 264744 334750
rect 264900 329118 264928 337742
rect 265084 335442 265112 337742
rect 265176 336258 265204 337878
rect 265164 336252 265216 336258
rect 265164 336194 265216 336200
rect 265268 336054 265296 338014
rect 265406 337770 265434 338028
rect 265498 337906 265526 338028
rect 265636 338014 265696 338042
rect 265498 337878 265572 337906
rect 265406 337742 265480 337770
rect 265452 336462 265480 337742
rect 265440 336456 265492 336462
rect 265440 336398 265492 336404
rect 265256 336048 265308 336054
rect 265256 335990 265308 335996
rect 265072 335436 265124 335442
rect 265072 335378 265124 335384
rect 265544 333266 265572 337878
rect 265636 333674 265664 338014
rect 265774 337770 265802 338028
rect 265866 337872 265894 338028
rect 266004 338014 266064 338042
rect 265866 337844 265940 337872
rect 265774 337742 265848 337770
rect 265820 336530 265848 337742
rect 265808 336524 265860 336530
rect 265808 336466 265860 336472
rect 265808 335436 265860 335442
rect 265808 335378 265860 335384
rect 265624 333668 265676 333674
rect 265624 333610 265676 333616
rect 265532 333260 265584 333266
rect 265532 333202 265584 333208
rect 264888 329112 264940 329118
rect 264888 329054 264940 329060
rect 264704 5024 264756 5030
rect 264704 4966 264756 4972
rect 265820 4826 265848 335378
rect 265912 328454 265940 337844
rect 266004 333538 266032 338014
rect 266142 337906 266170 338028
rect 266096 337878 266170 337906
rect 266096 335986 266124 337878
rect 266234 337770 266262 338028
rect 266188 337742 266262 337770
rect 266372 338014 266432 338042
rect 266084 335980 266136 335986
rect 266084 335922 266136 335928
rect 265992 333532 266044 333538
rect 265992 333474 266044 333480
rect 266084 333260 266136 333266
rect 266084 333202 266136 333208
rect 265912 328426 266032 328454
rect 265900 328296 265952 328302
rect 265900 328238 265952 328244
rect 265912 9246 265940 328238
rect 266004 9314 266032 328426
rect 266096 9382 266124 333202
rect 266188 328302 266216 337742
rect 266372 331430 266400 338014
rect 266510 337770 266538 338028
rect 266602 337872 266630 338028
rect 266740 338014 266800 338042
rect 266602 337844 266676 337872
rect 266510 337742 266584 337770
rect 266556 336598 266584 337742
rect 266544 336592 266596 336598
rect 266544 336534 266596 336540
rect 266648 335492 266676 337844
rect 266740 335646 266768 338014
rect 266878 337770 266906 338028
rect 266970 337872 266998 338028
rect 267108 338014 267168 338042
rect 266970 337844 267044 337872
rect 266878 337742 266952 337770
rect 266924 336326 266952 337742
rect 266912 336320 266964 336326
rect 266912 336262 266964 336268
rect 267016 336172 267044 337844
rect 266924 336144 267044 336172
rect 266728 335640 266780 335646
rect 266728 335582 266780 335588
rect 266648 335464 266768 335492
rect 266636 335368 266688 335374
rect 266636 335310 266688 335316
rect 266360 331424 266412 331430
rect 266360 331366 266412 331372
rect 266176 328296 266228 328302
rect 266176 328238 266228 328244
rect 266648 325446 266676 335310
rect 266740 332722 266768 335464
rect 266924 332790 266952 336144
rect 267004 335912 267056 335918
rect 267004 335854 267056 335860
rect 266912 332784 266964 332790
rect 266912 332726 266964 332732
rect 266728 332716 266780 332722
rect 266728 332658 266780 332664
rect 266636 325440 266688 325446
rect 266636 325382 266688 325388
rect 266084 9376 266136 9382
rect 266084 9318 266136 9324
rect 265992 9308 266044 9314
rect 265992 9250 266044 9256
rect 265900 9240 265952 9246
rect 265900 9182 265952 9188
rect 267016 6186 267044 335854
rect 267108 335374 267136 338014
rect 267246 337770 267274 338028
rect 267338 337872 267366 338028
rect 267476 338014 267536 338042
rect 267338 337844 267412 337872
rect 267200 337742 267274 337770
rect 267096 335368 267148 335374
rect 267096 335310 267148 335316
rect 267200 334218 267228 337742
rect 267280 335368 267332 335374
rect 267280 335310 267332 335316
rect 267188 334212 267240 334218
rect 267188 334154 267240 334160
rect 267188 330540 267240 330546
rect 267188 330482 267240 330488
rect 267200 15910 267228 330482
rect 267188 15904 267240 15910
rect 267188 15846 267240 15852
rect 267004 6180 267056 6186
rect 267004 6122 267056 6128
rect 267292 4962 267320 335310
rect 267384 331498 267412 337844
rect 267372 331492 267424 331498
rect 267372 331434 267424 331440
rect 267476 330546 267504 338014
rect 267614 337906 267642 338028
rect 267568 337878 267642 337906
rect 267568 334286 267596 337878
rect 267706 337770 267734 338028
rect 267660 337742 267734 337770
rect 267844 338014 267904 338042
rect 267556 334280 267608 334286
rect 267556 334222 267608 334228
rect 267464 330540 267516 330546
rect 267464 330482 267516 330488
rect 267660 330274 267688 337742
rect 267844 335374 267872 338014
rect 267982 337770 268010 338028
rect 268074 337872 268102 338028
rect 268212 338014 268272 338042
rect 268074 337844 268148 337872
rect 267982 337742 268056 337770
rect 268028 335578 268056 337742
rect 268016 335572 268068 335578
rect 268016 335514 268068 335520
rect 267832 335368 267884 335374
rect 267832 335310 267884 335316
rect 268120 332858 268148 337844
rect 268212 335374 268240 338014
rect 268350 337770 268378 338028
rect 268442 337872 268470 338028
rect 268580 338014 268640 338042
rect 268442 337844 268516 337872
rect 268350 337742 268424 337770
rect 268200 335368 268252 335374
rect 268200 335310 268252 335316
rect 268396 334354 268424 337742
rect 268384 334348 268436 334354
rect 268384 334290 268436 334296
rect 268108 332852 268160 332858
rect 268108 332794 268160 332800
rect 268488 331566 268516 337844
rect 268476 331560 268528 331566
rect 268476 331502 268528 331508
rect 267648 330268 267700 330274
rect 267648 330210 267700 330216
rect 268580 316034 268608 338014
rect 268718 337906 268746 338028
rect 268672 337878 268746 337906
rect 268672 336190 268700 337878
rect 268810 337770 268838 338028
rect 268902 337906 268930 338028
rect 269040 338014 269100 338042
rect 268902 337878 268976 337906
rect 268764 337742 268838 337770
rect 268660 336184 268712 336190
rect 268660 336126 268712 336132
rect 268660 335436 268712 335442
rect 268660 335378 268712 335384
rect 268488 316006 268608 316034
rect 268488 9178 268516 316006
rect 268476 9172 268528 9178
rect 268476 9114 268528 9120
rect 268672 5710 268700 335378
rect 268764 335374 268792 337742
rect 268948 335458 268976 337878
rect 268856 335430 268976 335458
rect 269040 335442 269068 338014
rect 269178 337770 269206 338028
rect 269270 337872 269298 338028
rect 269270 337844 269344 337872
rect 269178 337742 269252 337770
rect 269028 335436 269080 335442
rect 268752 335368 268804 335374
rect 268752 335310 268804 335316
rect 268752 335232 268804 335238
rect 268752 335174 268804 335180
rect 268764 325378 268792 335174
rect 268752 325372 268804 325378
rect 268752 325314 268804 325320
rect 268856 323950 268884 335430
rect 269028 335378 269080 335384
rect 268936 335368 268988 335374
rect 268936 335310 268988 335316
rect 268948 330342 268976 335310
rect 269224 334422 269252 337742
rect 269212 334416 269264 334422
rect 269212 334358 269264 334364
rect 269316 332926 269344 337844
rect 269454 337770 269482 338028
rect 269546 337872 269574 338028
rect 269638 337940 269666 338028
rect 269638 337912 269712 337940
rect 269546 337844 269620 337872
rect 269454 337742 269528 337770
rect 269304 332920 269356 332926
rect 269304 332862 269356 332868
rect 268936 330336 268988 330342
rect 268936 330278 268988 330284
rect 269500 325694 269528 337742
rect 269592 335714 269620 337844
rect 269580 335708 269632 335714
rect 269580 335650 269632 335656
rect 269684 331702 269712 337912
rect 269822 337770 269850 338028
rect 269914 337890 269942 338028
rect 270006 337940 270034 338028
rect 270144 338014 270204 338042
rect 270006 337912 270080 337940
rect 269902 337884 269954 337890
rect 269902 337826 269954 337832
rect 269822 337742 269896 337770
rect 269764 335504 269816 335510
rect 269764 335446 269816 335452
rect 269672 331696 269724 331702
rect 269672 331638 269724 331644
rect 269776 325694 269804 335446
rect 269868 330562 269896 337742
rect 269868 330534 269988 330562
rect 269500 325666 269712 325694
rect 269776 325666 269896 325694
rect 268844 323944 268896 323950
rect 268844 323886 268896 323892
rect 269684 5778 269712 325666
rect 269868 5914 269896 325666
rect 269856 5908 269908 5914
rect 269856 5850 269908 5856
rect 269960 5846 269988 330534
rect 270052 328982 270080 337912
rect 270144 335510 270172 338014
rect 270282 337770 270310 338028
rect 270374 337906 270402 338028
rect 270374 337878 270448 337906
rect 270236 337742 270310 337770
rect 270132 335504 270184 335510
rect 270132 335446 270184 335452
rect 270040 328976 270092 328982
rect 270040 328918 270092 328924
rect 270236 328794 270264 337742
rect 270420 330410 270448 337878
rect 270558 337770 270586 338028
rect 270650 337890 270678 338028
rect 270742 337906 270770 338028
rect 270880 338014 270940 338042
rect 270638 337884 270690 337890
rect 270742 337878 270816 337906
rect 270638 337826 270690 337832
rect 270558 337742 270632 337770
rect 270500 335368 270552 335374
rect 270500 335310 270552 335316
rect 270408 330404 270460 330410
rect 270408 330346 270460 330352
rect 270052 328766 270264 328794
rect 270052 9858 270080 328766
rect 270132 328704 270184 328710
rect 270132 328646 270184 328652
rect 270040 9852 270092 9858
rect 270040 9794 270092 9800
rect 270144 9790 270172 328646
rect 270512 325694 270540 335310
rect 270604 331214 270632 337742
rect 270788 337686 270816 337878
rect 270776 337680 270828 337686
rect 270776 337622 270828 337628
rect 270880 334370 270908 338014
rect 271018 337770 271046 338028
rect 270972 337742 271046 337770
rect 270972 335374 271000 337742
rect 271110 337634 271138 338028
rect 271064 337606 271138 337634
rect 271248 338014 271308 338042
rect 270960 335368 271012 335374
rect 270960 335310 271012 335316
rect 271064 334490 271092 337606
rect 271248 335374 271276 338014
rect 271386 337770 271414 338028
rect 271478 337890 271506 338028
rect 271616 338014 271676 338042
rect 271466 337884 271518 337890
rect 271466 337826 271518 337832
rect 271386 337742 271460 337770
rect 271328 335436 271380 335442
rect 271328 335378 271380 335384
rect 271236 335368 271288 335374
rect 271236 335310 271288 335316
rect 271340 334642 271368 335378
rect 271156 334614 271368 334642
rect 271052 334484 271104 334490
rect 271052 334426 271104 334432
rect 270880 334342 271092 334370
rect 270604 331186 270908 331214
rect 270880 325694 270908 331186
rect 270512 325666 270632 325694
rect 270880 325666 271000 325694
rect 270604 9994 270632 325666
rect 270592 9988 270644 9994
rect 270592 9930 270644 9936
rect 270132 9784 270184 9790
rect 270132 9726 270184 9732
rect 270972 5982 271000 325666
rect 271064 6050 271092 334342
rect 271156 10130 271184 334614
rect 271328 334552 271380 334558
rect 271328 334494 271380 334500
rect 271144 10124 271196 10130
rect 271144 10066 271196 10072
rect 271340 9926 271368 334494
rect 271432 10062 271460 337742
rect 271512 335368 271564 335374
rect 271512 335310 271564 335316
rect 271420 10056 271472 10062
rect 271420 9998 271472 10004
rect 271328 9920 271380 9926
rect 271328 9862 271380 9868
rect 271524 6118 271552 335310
rect 271616 6730 271644 338014
rect 271754 337770 271782 338028
rect 271708 337742 271782 337770
rect 271708 335442 271736 337742
rect 271846 337634 271874 338028
rect 271800 337606 271874 337634
rect 271984 338014 272044 338042
rect 271800 335594 271828 337606
rect 271800 335566 271920 335594
rect 271696 335436 271748 335442
rect 271696 335378 271748 335384
rect 271892 335374 271920 335566
rect 271984 335510 272012 338014
rect 272122 337770 272150 338028
rect 272214 337906 272242 338028
rect 272352 338014 272412 338042
rect 272214 337878 272288 337906
rect 272122 337742 272196 337770
rect 271972 335504 272024 335510
rect 271972 335446 272024 335452
rect 271880 335368 271932 335374
rect 271880 335310 271932 335316
rect 271696 335300 271748 335306
rect 271696 335242 271748 335248
rect 271708 331770 271736 335242
rect 271696 331764 271748 331770
rect 271696 331706 271748 331712
rect 272168 330478 272196 337742
rect 272260 337618 272288 337878
rect 272248 337612 272300 337618
rect 272248 337554 272300 337560
rect 272352 335442 272380 338014
rect 272490 337770 272518 338028
rect 272582 337890 272610 338028
rect 272674 337906 272702 338028
rect 272812 338014 272872 338042
rect 272570 337884 272622 337890
rect 272674 337878 272748 337906
rect 272570 337826 272622 337832
rect 272490 337742 272564 337770
rect 272340 335436 272392 335442
rect 272340 335378 272392 335384
rect 272156 330472 272208 330478
rect 272156 330414 272208 330420
rect 272536 10266 272564 337742
rect 272616 336660 272668 336666
rect 272616 336602 272668 336608
rect 272628 10946 272656 336602
rect 272720 333266 272748 337878
rect 272708 333260 272760 333266
rect 272708 333202 272760 333208
rect 272812 330562 272840 338014
rect 272950 337906 272978 338028
rect 272904 337878 272978 337906
rect 272904 337482 272932 337878
rect 273042 337770 273070 338028
rect 272996 337742 273070 337770
rect 273180 338014 273240 338042
rect 272892 337476 272944 337482
rect 272892 337418 272944 337424
rect 272892 336048 272944 336054
rect 272890 336016 272892 336025
rect 272944 336016 272946 336025
rect 272890 335951 272946 335960
rect 272892 335844 272944 335850
rect 272892 335786 272944 335792
rect 272904 335617 272932 335786
rect 272890 335608 272946 335617
rect 272890 335543 272946 335552
rect 272892 335504 272944 335510
rect 272892 335446 272944 335452
rect 272904 330818 272932 335446
rect 272892 330812 272944 330818
rect 272892 330754 272944 330760
rect 272996 330698 273024 337742
rect 273180 336666 273208 338014
rect 273318 337906 273346 338028
rect 273272 337878 273346 337906
rect 273168 336660 273220 336666
rect 273168 336602 273220 336608
rect 273076 335436 273128 335442
rect 273076 335378 273128 335384
rect 272720 330534 272840 330562
rect 272904 330670 273024 330698
rect 272720 11014 272748 330534
rect 272800 330472 272852 330478
rect 272800 330414 272852 330420
rect 272708 11008 272760 11014
rect 272708 10950 272760 10956
rect 272616 10940 272668 10946
rect 272616 10882 272668 10888
rect 272524 10260 272576 10266
rect 272524 10202 272576 10208
rect 272812 10198 272840 330414
rect 272800 10192 272852 10198
rect 272800 10134 272852 10140
rect 271604 6724 271656 6730
rect 271604 6666 271656 6672
rect 272904 6458 272932 330670
rect 273088 330562 273116 335378
rect 273272 334694 273300 337878
rect 273410 337770 273438 338028
rect 273364 337742 273438 337770
rect 273548 338014 273608 338042
rect 273364 335510 273392 337742
rect 273444 337544 273496 337550
rect 273444 337486 273496 337492
rect 273352 335504 273404 335510
rect 273352 335446 273404 335452
rect 273260 334688 273312 334694
rect 273260 334630 273312 334636
rect 273168 333260 273220 333266
rect 273168 333202 273220 333208
rect 272996 330534 273116 330562
rect 272996 6594 273024 330534
rect 273076 330472 273128 330478
rect 273076 330414 273128 330420
rect 273088 6662 273116 330414
rect 273076 6656 273128 6662
rect 273076 6598 273128 6604
rect 272984 6588 273036 6594
rect 272984 6530 273036 6536
rect 273180 6526 273208 333202
rect 273456 328438 273484 337486
rect 273444 328432 273496 328438
rect 273444 328374 273496 328380
rect 273548 326398 273576 338014
rect 273686 337906 273714 338028
rect 273640 337878 273714 337906
rect 273640 335374 273668 337878
rect 273778 337770 273806 338028
rect 273732 337742 273806 337770
rect 273916 338014 273976 338042
rect 273628 335368 273680 335374
rect 273628 335310 273680 335316
rect 273628 334620 273680 334626
rect 273628 334562 273680 334568
rect 273640 329050 273668 334562
rect 273628 329044 273680 329050
rect 273628 328986 273680 328992
rect 273536 326392 273588 326398
rect 273536 326334 273588 326340
rect 273168 6520 273220 6526
rect 273168 6462 273220 6468
rect 272892 6452 272944 6458
rect 272892 6394 272944 6400
rect 273732 6322 273760 337742
rect 273916 336410 273944 338014
rect 274054 337634 274082 338028
rect 274146 337906 274174 338028
rect 274284 338014 274344 338042
rect 274146 337878 274220 337906
rect 273824 336382 273944 336410
rect 274008 337606 274082 337634
rect 273824 336326 273852 336382
rect 273812 336320 273864 336326
rect 273812 336262 273864 336268
rect 274008 334626 274036 337606
rect 274088 335368 274140 335374
rect 274088 335310 274140 335316
rect 273996 334620 274048 334626
rect 273996 334562 274048 334568
rect 273904 333260 273956 333266
rect 273904 333202 273956 333208
rect 273812 326460 273864 326466
rect 273812 326402 273864 326408
rect 273720 6316 273772 6322
rect 273720 6258 273772 6264
rect 273824 6186 273852 326402
rect 273916 6254 273944 333202
rect 274100 330478 274128 335310
rect 274192 333266 274220 337878
rect 274180 333260 274232 333266
rect 274180 333202 274232 333208
rect 274284 331214 274312 338014
rect 274422 337958 274450 338028
rect 274410 337952 274462 337958
rect 274410 337894 274462 337900
rect 274514 337906 274542 338028
rect 274652 338014 274712 338042
rect 274514 337878 274588 337906
rect 274364 336320 274416 336326
rect 274364 336262 274416 336268
rect 274192 331186 274312 331214
rect 274088 330472 274140 330478
rect 274088 330414 274140 330420
rect 273996 326392 274048 326398
rect 274192 326346 274220 331186
rect 273996 326334 274048 326340
rect 274008 10878 274036 326334
rect 274100 326318 274220 326346
rect 273996 10872 274048 10878
rect 273996 10814 274048 10820
rect 274100 10742 274128 326318
rect 274376 321554 274404 336262
rect 274456 335300 274508 335306
rect 274456 335242 274508 335248
rect 274192 321526 274404 321554
rect 274192 10810 274220 321526
rect 274468 316034 274496 335242
rect 274560 326466 274588 337878
rect 274652 335374 274680 338014
rect 274790 337770 274818 338028
rect 274882 337906 274910 338028
rect 275020 338014 275080 338042
rect 274882 337878 274956 337906
rect 274790 337742 274864 337770
rect 274640 335368 274692 335374
rect 274640 335310 274692 335316
rect 274836 331838 274864 337742
rect 274928 336161 274956 337878
rect 274914 336152 274970 336161
rect 274914 336087 274970 336096
rect 274824 331832 274876 331838
rect 274824 331774 274876 331780
rect 274548 326460 274600 326466
rect 274548 326402 274600 326408
rect 275020 326398 275048 338014
rect 275158 337906 275186 338028
rect 275112 337878 275186 337906
rect 275112 329798 275140 337878
rect 275250 337770 275278 338028
rect 275204 337742 275278 337770
rect 275388 338014 275448 338042
rect 275204 335442 275232 337742
rect 275282 337648 275338 337657
rect 275282 337583 275338 337592
rect 275192 335436 275244 335442
rect 275192 335378 275244 335384
rect 275296 331214 275324 337583
rect 275388 335458 275416 338014
rect 275526 337770 275554 338028
rect 275618 337906 275646 338028
rect 275756 338014 275816 338042
rect 275756 337929 275784 338014
rect 275742 337920 275798 337929
rect 275618 337878 275692 337906
rect 275526 337742 275600 337770
rect 275572 335594 275600 337742
rect 275664 335753 275692 337878
rect 275742 337855 275798 337864
rect 275894 337770 275922 338028
rect 275848 337742 275922 337770
rect 275650 335744 275706 335753
rect 275650 335679 275706 335688
rect 275572 335566 275784 335594
rect 275388 335430 275692 335458
rect 275468 335368 275520 335374
rect 275468 335310 275520 335316
rect 275204 331186 275324 331214
rect 275100 329792 275152 329798
rect 275100 329734 275152 329740
rect 275008 326392 275060 326398
rect 275008 326334 275060 326340
rect 275204 321554 275232 331186
rect 275376 326392 275428 326398
rect 275376 326334 275428 326340
rect 275204 321526 275324 321554
rect 274284 316006 274496 316034
rect 274180 10804 274232 10810
rect 274180 10746 274232 10752
rect 274088 10736 274140 10742
rect 274088 10678 274140 10684
rect 274284 6390 274312 316006
rect 275296 10470 275324 321526
rect 275388 10606 275416 326334
rect 275480 10674 275508 335310
rect 275560 334552 275612 334558
rect 275560 334494 275612 334500
rect 275572 326942 275600 334494
rect 275560 326936 275612 326942
rect 275560 326878 275612 326884
rect 275468 10668 275520 10674
rect 275468 10610 275520 10616
rect 275376 10600 275428 10606
rect 275376 10542 275428 10548
rect 275664 10538 275692 335430
rect 275756 328370 275784 335566
rect 275848 334558 275876 337742
rect 275986 337634 276014 338028
rect 275940 337606 276014 337634
rect 276124 338014 276184 338042
rect 275940 335374 275968 337606
rect 275928 335368 275980 335374
rect 275928 335310 275980 335316
rect 275836 334552 275888 334558
rect 275836 334494 275888 334500
rect 275744 328364 275796 328370
rect 275744 328306 275796 328312
rect 276124 321554 276152 338014
rect 276262 337770 276290 338028
rect 276354 337958 276382 338028
rect 276342 337952 276394 337958
rect 276342 337894 276394 337900
rect 276446 337906 276474 338028
rect 276446 337878 276520 337906
rect 276262 337742 276336 337770
rect 276308 325310 276336 337742
rect 276492 333266 276520 337878
rect 276630 337770 276658 338028
rect 276722 337958 276750 338028
rect 276710 337952 276762 337958
rect 276710 337894 276762 337900
rect 276814 337906 276842 338028
rect 276814 337878 276888 337906
rect 276630 337742 276704 337770
rect 276480 333260 276532 333266
rect 276480 333202 276532 333208
rect 276296 325304 276348 325310
rect 276296 325246 276348 325252
rect 276676 323882 276704 337742
rect 276756 335436 276808 335442
rect 276756 335378 276808 335384
rect 276664 323876 276716 323882
rect 276664 323818 276716 323824
rect 276124 321526 276612 321554
rect 275652 10532 275704 10538
rect 275652 10474 275704 10480
rect 275284 10464 275336 10470
rect 275284 10406 275336 10412
rect 276584 10402 276612 321526
rect 276572 10396 276624 10402
rect 276572 10338 276624 10344
rect 274272 6384 274324 6390
rect 274272 6326 274324 6332
rect 273904 6248 273956 6254
rect 273904 6190 273956 6196
rect 273628 6180 273680 6186
rect 273628 6122 273680 6128
rect 273812 6180 273864 6186
rect 273812 6122 273864 6128
rect 271512 6112 271564 6118
rect 271512 6054 271564 6060
rect 271052 6044 271104 6050
rect 271052 5986 271104 5992
rect 270960 5976 271012 5982
rect 270960 5918 271012 5924
rect 269948 5840 270000 5846
rect 269948 5782 270000 5788
rect 269672 5772 269724 5778
rect 269672 5714 269724 5720
rect 268660 5704 268712 5710
rect 268660 5646 268712 5652
rect 267740 5500 267792 5506
rect 267740 5442 267792 5448
rect 272432 5500 272484 5506
rect 272432 5442 272484 5448
rect 267280 4956 267332 4962
rect 267280 4898 267332 4904
rect 265808 4820 265860 4826
rect 265808 4762 265860 4768
rect 266544 3596 266596 3602
rect 266544 3538 266596 3544
rect 264244 3528 264296 3534
rect 264244 3470 264296 3476
rect 265348 3528 265400 3534
rect 265348 3470 265400 3476
rect 264152 3460 264204 3466
rect 264152 3402 264204 3408
rect 263508 3188 263560 3194
rect 263508 3130 263560 3136
rect 263324 3052 263376 3058
rect 263324 2994 263376 3000
rect 264164 480 264192 3402
rect 265360 480 265388 3470
rect 266556 480 266584 3538
rect 267752 480 267780 5442
rect 271236 4684 271288 4690
rect 271236 4626 271288 4632
rect 270040 3188 270092 3194
rect 270040 3130 270092 3136
rect 268844 3052 268896 3058
rect 268844 2994 268896 3000
rect 268856 480 268884 2994
rect 270052 480 270080 3130
rect 271248 480 271276 4626
rect 272444 480 272472 5442
rect 273640 480 273668 6122
rect 276020 5432 276072 5438
rect 276020 5374 276072 5380
rect 274824 4752 274876 4758
rect 274824 4694 274876 4700
rect 274836 480 274864 4694
rect 276032 480 276060 5374
rect 276768 2922 276796 335378
rect 276860 329730 276888 337878
rect 276998 337770 277026 338028
rect 277090 337958 277118 338028
rect 277078 337952 277130 337958
rect 277078 337894 277130 337900
rect 277182 337906 277210 338028
rect 277320 338014 277380 338042
rect 277182 337878 277256 337906
rect 276998 337742 277072 337770
rect 276940 335776 276992 335782
rect 276940 335718 276992 335724
rect 276952 331634 276980 335718
rect 276940 331628 276992 331634
rect 276940 331570 276992 331576
rect 276848 329724 276900 329730
rect 276848 329666 276900 329672
rect 277044 322386 277072 337742
rect 277124 333260 277176 333266
rect 277124 333202 277176 333208
rect 277032 322380 277084 322386
rect 277032 322322 277084 322328
rect 277136 10334 277164 333202
rect 277228 329662 277256 337878
rect 277320 335442 277348 338014
rect 277458 337770 277486 338028
rect 277550 337872 277578 338028
rect 277688 338014 277748 338042
rect 277550 337844 277624 337872
rect 277412 337742 277486 337770
rect 277412 336326 277440 337742
rect 277492 336388 277544 336394
rect 277492 336330 277544 336336
rect 277400 336320 277452 336326
rect 277400 336262 277452 336268
rect 277308 335436 277360 335442
rect 277308 335378 277360 335384
rect 277504 331214 277532 336330
rect 277596 333266 277624 337844
rect 277688 335510 277716 338014
rect 277826 337906 277854 338028
rect 277780 337878 277854 337906
rect 277676 335504 277728 335510
rect 277676 335446 277728 335452
rect 277780 335170 277808 337878
rect 277918 337770 277946 338028
rect 277872 337742 277946 337770
rect 278102 337770 278130 338028
rect 278194 337890 278222 338028
rect 278182 337884 278234 337890
rect 278182 337826 278234 337832
rect 278286 337770 278314 338028
rect 278102 337742 278176 337770
rect 277768 335164 277820 335170
rect 277768 335106 277820 335112
rect 277584 333260 277636 333266
rect 277584 333202 277636 333208
rect 277504 331186 277716 331214
rect 277216 329656 277268 329662
rect 277216 329598 277268 329604
rect 277124 10328 277176 10334
rect 277124 10270 277176 10276
rect 277688 4418 277716 331186
rect 277872 328234 277900 337742
rect 278148 335492 278176 337742
rect 278056 335464 278176 335492
rect 278240 337742 278314 337770
rect 278424 338014 278484 338042
rect 277860 328228 277912 328234
rect 277860 328170 277912 328176
rect 278056 316034 278084 335464
rect 278136 335368 278188 335374
rect 278136 335310 278188 335316
rect 277964 316006 278084 316034
rect 277124 4412 277176 4418
rect 277124 4354 277176 4360
rect 277676 4412 277728 4418
rect 277676 4354 277728 4360
rect 276756 2916 276808 2922
rect 276756 2858 276808 2864
rect 277136 480 277164 4354
rect 277964 3058 277992 316006
rect 278148 3126 278176 335310
rect 278240 328166 278268 337742
rect 278318 336016 278374 336025
rect 278318 335951 278374 335960
rect 278332 335782 278360 335951
rect 278320 335776 278372 335782
rect 278320 335718 278372 335724
rect 278318 335608 278374 335617
rect 278318 335543 278320 335552
rect 278372 335543 278374 335552
rect 278320 335514 278372 335520
rect 278424 335374 278452 338014
rect 278562 337906 278590 338028
rect 278516 337878 278590 337906
rect 278516 335714 278544 337878
rect 278654 337770 278682 338028
rect 278608 337742 278682 337770
rect 278792 338014 278852 338042
rect 278504 335708 278556 335714
rect 278504 335650 278556 335656
rect 278504 335504 278556 335510
rect 278504 335446 278556 335452
rect 278412 335368 278464 335374
rect 278412 335310 278464 335316
rect 278320 333260 278372 333266
rect 278320 333202 278372 333208
rect 278332 328302 278360 333202
rect 278320 328296 278372 328302
rect 278320 328238 278372 328244
rect 278228 328160 278280 328166
rect 278228 328102 278280 328108
rect 278320 5364 278372 5370
rect 278320 5306 278372 5312
rect 278136 3120 278188 3126
rect 278136 3062 278188 3068
rect 277952 3052 278004 3058
rect 277952 2994 278004 3000
rect 278332 480 278360 5306
rect 278516 2990 278544 335446
rect 278608 326874 278636 337742
rect 278688 335708 278740 335714
rect 278688 335650 278740 335656
rect 278700 333878 278728 335650
rect 278792 335374 278820 338014
rect 278930 337770 278958 338028
rect 279022 337906 279050 338028
rect 279160 338014 279220 338042
rect 279022 337878 279096 337906
rect 278930 337742 279004 337770
rect 278976 337414 279004 337742
rect 278964 337408 279016 337414
rect 278964 337350 279016 337356
rect 279068 337346 279096 337878
rect 279056 337340 279108 337346
rect 279056 337282 279108 337288
rect 279160 335442 279188 338014
rect 279298 337770 279326 338028
rect 279390 337906 279418 338028
rect 279528 338014 279588 338042
rect 279390 337878 279464 337906
rect 279298 337742 279372 337770
rect 279344 335617 279372 337742
rect 279436 337278 279464 337878
rect 279424 337272 279476 337278
rect 279424 337214 279476 337220
rect 279528 335714 279556 338014
rect 279666 337770 279694 338028
rect 279758 337906 279786 338028
rect 279758 337878 279832 337906
rect 279620 337742 279694 337770
rect 279516 335708 279568 335714
rect 279516 335650 279568 335656
rect 279330 335608 279386 335617
rect 279330 335543 279386 335552
rect 279148 335436 279200 335442
rect 279148 335378 279200 335384
rect 278780 335368 278832 335374
rect 278780 335310 278832 335316
rect 279516 335368 279568 335374
rect 279516 335310 279568 335316
rect 278688 333872 278740 333878
rect 278688 333814 278740 333820
rect 278596 326868 278648 326874
rect 278596 326810 278648 326816
rect 279528 321554 279556 335310
rect 279620 335102 279648 337742
rect 279700 335708 279752 335714
rect 279700 335650 279752 335656
rect 279608 335096 279660 335102
rect 279608 335038 279660 335044
rect 279712 321554 279740 335650
rect 279804 331226 279832 337878
rect 279942 337770 279970 338028
rect 280034 337890 280062 338028
rect 280022 337884 280074 337890
rect 280022 337826 280074 337832
rect 280126 337770 280154 338028
rect 280218 337906 280246 338028
rect 280356 338014 280416 338042
rect 280218 337878 280292 337906
rect 279942 337742 280016 337770
rect 279884 335436 279936 335442
rect 279884 335378 279936 335384
rect 279792 331220 279844 331226
rect 279792 331162 279844 331168
rect 279528 321526 279648 321554
rect 279712 321526 279832 321554
rect 279516 5296 279568 5302
rect 279516 5238 279568 5244
rect 278504 2984 278556 2990
rect 278504 2926 278556 2932
rect 279528 480 279556 5238
rect 279620 3194 279648 321526
rect 279804 3330 279832 321526
rect 279792 3324 279844 3330
rect 279792 3266 279844 3272
rect 279896 3262 279924 335378
rect 279988 3398 280016 337742
rect 280080 337742 280154 337770
rect 280080 329594 280108 337742
rect 280264 333266 280292 337878
rect 280252 333260 280304 333266
rect 280252 333202 280304 333208
rect 280068 329588 280120 329594
rect 280068 329530 280120 329536
rect 280356 326398 280384 338014
rect 280494 337770 280522 338028
rect 280586 337906 280614 338028
rect 280724 338014 280784 338042
rect 280586 337878 280660 337906
rect 280494 337742 280568 337770
rect 280436 337204 280488 337210
rect 280436 337146 280488 337152
rect 280344 326392 280396 326398
rect 280344 326334 280396 326340
rect 280448 321554 280476 337146
rect 280540 326482 280568 337742
rect 280632 333334 280660 337878
rect 280724 336802 280752 338014
rect 280862 337770 280890 338028
rect 280954 337822 280982 338028
rect 281092 338014 281152 338042
rect 280816 337742 280890 337770
rect 280942 337816 280994 337822
rect 280942 337758 280994 337764
rect 280712 336796 280764 336802
rect 280712 336738 280764 336744
rect 280816 335594 280844 337742
rect 280896 336796 280948 336802
rect 280896 336738 280948 336744
rect 280724 335566 280844 335594
rect 280620 333328 280672 333334
rect 280620 333270 280672 333276
rect 280724 331214 280752 335566
rect 280804 335436 280856 335442
rect 280804 335378 280856 335384
rect 280632 331186 280752 331214
rect 280632 326602 280660 331186
rect 280620 326596 280672 326602
rect 280620 326538 280672 326544
rect 280540 326454 280752 326482
rect 280620 326324 280672 326330
rect 280620 326266 280672 326272
rect 280448 321526 280568 321554
rect 280540 12034 280568 321526
rect 280632 12102 280660 326266
rect 280724 12170 280752 326454
rect 280712 12164 280764 12170
rect 280712 12106 280764 12112
rect 280620 12096 280672 12102
rect 280620 12038 280672 12044
rect 280528 12028 280580 12034
rect 280528 11970 280580 11976
rect 280816 7818 280844 335378
rect 280908 7954 280936 336738
rect 280988 326392 281040 326398
rect 280988 326334 281040 326340
rect 281000 8022 281028 326334
rect 280988 8016 281040 8022
rect 280988 7958 281040 7964
rect 280896 7948 280948 7954
rect 280896 7890 280948 7896
rect 281092 7886 281120 338014
rect 281230 337958 281258 338028
rect 281218 337952 281270 337958
rect 281322 337940 281350 338028
rect 281460 338014 281520 338042
rect 281322 337912 281396 337940
rect 281218 337894 281270 337900
rect 281172 337816 281224 337822
rect 281172 337758 281224 337764
rect 281080 7880 281132 7886
rect 281080 7822 281132 7828
rect 280804 7812 280856 7818
rect 280804 7754 280856 7760
rect 280712 4208 280764 4214
rect 280712 4150 280764 4156
rect 279976 3392 280028 3398
rect 279976 3334 280028 3340
rect 279884 3256 279936 3262
rect 279884 3198 279936 3204
rect 279608 3188 279660 3194
rect 279608 3130 279660 3136
rect 280724 480 280752 4150
rect 281184 4010 281212 337758
rect 281264 333328 281316 333334
rect 281264 333270 281316 333276
rect 281276 4078 281304 333270
rect 281368 326466 281396 337912
rect 281460 335442 281488 338014
rect 281598 337770 281626 338028
rect 281690 337872 281718 338028
rect 281828 338014 281888 338042
rect 281690 337844 281764 337872
rect 281598 337742 281672 337770
rect 281448 335436 281500 335442
rect 281448 335378 281500 335384
rect 281448 333260 281500 333266
rect 281448 333202 281500 333208
rect 281356 326460 281408 326466
rect 281356 326402 281408 326408
rect 281460 326346 281488 333202
rect 281368 326318 281488 326346
rect 281368 4146 281396 326318
rect 281448 326256 281500 326262
rect 281448 326198 281500 326204
rect 281356 4140 281408 4146
rect 281356 4082 281408 4088
rect 281264 4072 281316 4078
rect 281264 4014 281316 4020
rect 281172 4004 281224 4010
rect 281172 3946 281224 3952
rect 281460 3942 281488 326198
rect 281644 321554 281672 337742
rect 281736 326194 281764 337844
rect 281724 326188 281776 326194
rect 281724 326130 281776 326136
rect 281828 326126 281856 338014
rect 281966 337906 281994 338028
rect 281920 337878 281994 337906
rect 282058 337906 282086 338028
rect 282196 338014 282256 338042
rect 282058 337878 282132 337906
rect 281920 331214 281948 337878
rect 282104 334762 282132 337878
rect 282196 335374 282224 338014
rect 282334 337906 282362 338028
rect 282288 337878 282362 337906
rect 282184 335368 282236 335374
rect 282184 335310 282236 335316
rect 282092 334756 282144 334762
rect 282092 334698 282144 334704
rect 282092 334620 282144 334626
rect 282092 334562 282144 334568
rect 281920 331186 282040 331214
rect 281816 326120 281868 326126
rect 281816 326062 281868 326068
rect 281644 321526 281948 321554
rect 281920 11966 281948 321526
rect 281908 11960 281960 11966
rect 281908 11902 281960 11908
rect 282012 11898 282040 331186
rect 282000 11892 282052 11898
rect 282000 11834 282052 11840
rect 282104 11762 282132 334562
rect 282288 331214 282316 337878
rect 282426 337770 282454 338028
rect 282564 338014 282624 338042
rect 282426 337742 282500 337770
rect 282472 335481 282500 337742
rect 282458 335472 282514 335481
rect 282458 335407 282514 335416
rect 282460 335368 282512 335374
rect 282460 335310 282512 335316
rect 282368 334756 282420 334762
rect 282368 334698 282420 334704
rect 282196 331186 282316 331214
rect 282196 11830 282224 331186
rect 282380 326618 282408 334698
rect 282288 326590 282408 326618
rect 282288 326262 282316 326590
rect 282368 326460 282420 326466
rect 282368 326402 282420 326408
rect 282276 326256 282328 326262
rect 282276 326198 282328 326204
rect 282276 326120 282328 326126
rect 282276 326062 282328 326068
rect 282184 11824 282236 11830
rect 282184 11766 282236 11772
rect 282092 11756 282144 11762
rect 282092 11698 282144 11704
rect 282288 7750 282316 326062
rect 282276 7744 282328 7750
rect 282276 7686 282328 7692
rect 282380 7614 282408 326402
rect 282472 7682 282500 335310
rect 282564 326466 282592 338014
rect 282702 337770 282730 338028
rect 282794 337906 282822 338028
rect 282932 338014 282992 338042
rect 282794 337878 282868 337906
rect 282702 337742 282776 337770
rect 282644 336456 282696 336462
rect 282644 336398 282696 336404
rect 282552 326460 282604 326466
rect 282552 326402 282604 326408
rect 282656 326346 282684 336398
rect 282748 334626 282776 337742
rect 282840 336462 282868 337878
rect 282828 336456 282880 336462
rect 282828 336398 282880 336404
rect 282826 336152 282882 336161
rect 282826 336087 282882 336096
rect 282840 335850 282868 336087
rect 282932 336025 282960 338014
rect 283070 337770 283098 338028
rect 283162 337906 283190 338028
rect 283300 338014 283360 338042
rect 283162 337878 283236 337906
rect 283070 337742 283144 337770
rect 282918 336016 282974 336025
rect 282918 335951 282974 335960
rect 282828 335844 282880 335850
rect 282828 335786 282880 335792
rect 282826 335744 282882 335753
rect 282826 335679 282882 335688
rect 282840 335646 282868 335679
rect 282828 335640 282880 335646
rect 282828 335582 282880 335588
rect 283116 335481 283144 337742
rect 282826 335472 282882 335481
rect 282826 335407 282882 335416
rect 283102 335472 283158 335481
rect 283102 335407 283158 335416
rect 282736 334620 282788 334626
rect 282736 334562 282788 334568
rect 282840 326346 282868 335407
rect 283208 333334 283236 337878
rect 283300 337142 283328 338014
rect 283438 337770 283466 338028
rect 283530 337906 283558 338028
rect 283668 338014 283728 338042
rect 283668 337958 283696 338014
rect 283656 337952 283708 337958
rect 283530 337878 283604 337906
rect 283656 337894 283708 337900
rect 283438 337742 283512 337770
rect 283288 337136 283340 337142
rect 283288 337078 283340 337084
rect 283484 337074 283512 337742
rect 283472 337068 283524 337074
rect 283472 337010 283524 337016
rect 283196 333328 283248 333334
rect 283196 333270 283248 333276
rect 283576 333266 283604 337878
rect 283806 337770 283834 338028
rect 283898 337804 283926 338028
rect 283990 337958 284018 338028
rect 284128 338014 284188 338042
rect 283978 337952 284030 337958
rect 283978 337894 284030 337900
rect 283898 337776 283972 337804
rect 283668 337742 283834 337770
rect 283564 333260 283616 333266
rect 283564 333202 283616 333208
rect 283668 329526 283696 337742
rect 283748 333328 283800 333334
rect 283748 333270 283800 333276
rect 283656 329520 283708 329526
rect 283656 329462 283708 329468
rect 282564 326318 282684 326346
rect 282748 326318 282868 326346
rect 282460 7676 282512 7682
rect 282460 7618 282512 7624
rect 282368 7608 282420 7614
rect 282368 7550 282420 7556
rect 281908 5228 281960 5234
rect 281908 5170 281960 5176
rect 281448 3936 281500 3942
rect 281448 3878 281500 3884
rect 281920 480 281948 5170
rect 282564 3670 282592 326318
rect 282644 326256 282696 326262
rect 282644 326198 282696 326204
rect 282656 3806 282684 326198
rect 282644 3800 282696 3806
rect 282644 3742 282696 3748
rect 282748 3738 282776 326318
rect 282828 326188 282880 326194
rect 282828 326130 282880 326136
rect 282840 3874 282868 326130
rect 283104 5160 283156 5166
rect 283104 5102 283156 5108
rect 282828 3868 282880 3874
rect 282828 3810 282880 3816
rect 282736 3732 282788 3738
rect 282736 3674 282788 3680
rect 282552 3664 282604 3670
rect 282552 3606 282604 3612
rect 283116 480 283144 5102
rect 283760 3602 283788 333270
rect 283944 331214 283972 337776
rect 284024 333260 284076 333266
rect 284024 333202 284076 333208
rect 283852 331186 283972 331214
rect 283852 326074 283880 331186
rect 284036 326346 284064 333202
rect 284128 327894 284156 338014
rect 284266 337770 284294 338028
rect 284358 337822 284386 338028
rect 284496 338014 284556 338042
rect 284220 337742 284294 337770
rect 284346 337816 284398 337822
rect 284346 337758 284398 337764
rect 284116 327888 284168 327894
rect 284116 327830 284168 327836
rect 284036 326318 284156 326346
rect 283852 326046 284064 326074
rect 283932 321632 283984 321638
rect 283932 321574 283984 321580
rect 283748 3596 283800 3602
rect 283748 3538 283800 3544
rect 283944 3534 283972 321574
rect 283932 3528 283984 3534
rect 283932 3470 283984 3476
rect 284036 3466 284064 326046
rect 284128 321638 284156 326318
rect 284116 321632 284168 321638
rect 284116 321574 284168 321580
rect 284220 316034 284248 337742
rect 284300 336116 284352 336122
rect 284300 336058 284352 336064
rect 284312 331214 284340 336058
rect 284496 335594 284524 338014
rect 284634 337770 284662 338028
rect 284726 337906 284754 338028
rect 284864 338014 284924 338042
rect 284726 337878 284800 337906
rect 284634 337742 284708 337770
rect 284496 335566 284616 335594
rect 284392 335504 284444 335510
rect 284392 335446 284444 335452
rect 284484 335504 284536 335510
rect 284484 335446 284536 335452
rect 284404 334762 284432 335446
rect 284392 334756 284444 334762
rect 284392 334698 284444 334704
rect 284312 331186 284432 331214
rect 284300 331016 284352 331022
rect 284300 330958 284352 330964
rect 284128 316006 284248 316034
rect 284128 3777 284156 316006
rect 284114 3768 284170 3777
rect 284114 3703 284170 3712
rect 284024 3460 284076 3466
rect 284024 3402 284076 3408
rect 284312 480 284340 330958
rect 284404 5506 284432 331186
rect 284496 9110 284524 335446
rect 284588 332450 284616 335566
rect 284680 335374 284708 337742
rect 284668 335368 284720 335374
rect 284668 335310 284720 335316
rect 284772 335034 284800 337878
rect 284864 336802 284892 338014
rect 285002 337770 285030 338028
rect 285094 337822 285122 338028
rect 284956 337742 285030 337770
rect 285082 337816 285134 337822
rect 285082 337758 285134 337764
rect 285278 337770 285306 338028
rect 285370 337872 285398 338028
rect 285462 337940 285490 338028
rect 285600 338014 285660 338042
rect 285462 337912 285536 337940
rect 285370 337844 285444 337872
rect 285278 337742 285352 337770
rect 284852 336796 284904 336802
rect 284852 336738 284904 336744
rect 284850 335608 284906 335617
rect 284850 335543 284906 335552
rect 284760 335028 284812 335034
rect 284760 334970 284812 334976
rect 284864 332586 284892 335543
rect 284852 332580 284904 332586
rect 284852 332522 284904 332528
rect 284576 332444 284628 332450
rect 284576 332386 284628 332392
rect 284956 326738 284984 337742
rect 285036 336796 285088 336802
rect 285036 336738 285088 336744
rect 285048 332382 285076 336738
rect 285128 336592 285180 336598
rect 285128 336534 285180 336540
rect 285140 334082 285168 336534
rect 285220 335776 285272 335782
rect 285220 335718 285272 335724
rect 285128 334076 285180 334082
rect 285128 334018 285180 334024
rect 285232 333062 285260 335718
rect 285220 333056 285272 333062
rect 285220 332998 285272 333004
rect 285036 332376 285088 332382
rect 285036 332318 285088 332324
rect 285324 331090 285352 337742
rect 285416 335510 285444 337844
rect 285508 335782 285536 337912
rect 285496 335776 285548 335782
rect 285496 335718 285548 335724
rect 285496 335572 285548 335578
rect 285496 335514 285548 335520
rect 285404 335504 285456 335510
rect 285404 335446 285456 335452
rect 285404 335368 285456 335374
rect 285404 335310 285456 335316
rect 285312 331084 285364 331090
rect 285312 331026 285364 331032
rect 285416 326806 285444 335310
rect 285508 334694 285536 335514
rect 285496 334688 285548 334694
rect 285496 334630 285548 334636
rect 285600 331022 285628 338014
rect 285738 337770 285766 338028
rect 285830 337906 285858 338028
rect 285968 338014 286028 338042
rect 285830 337878 285904 337906
rect 285738 337742 285812 337770
rect 285680 335436 285732 335442
rect 285680 335378 285732 335384
rect 285692 331214 285720 335378
rect 285784 335374 285812 337742
rect 285876 336666 285904 337878
rect 285864 336660 285916 336666
rect 285864 336602 285916 336608
rect 285968 336122 285996 338014
rect 286106 337770 286134 338028
rect 286198 337822 286226 338028
rect 286336 338014 286396 338042
rect 286060 337742 286134 337770
rect 286186 337816 286238 337822
rect 286186 337758 286238 337764
rect 285956 336116 286008 336122
rect 285956 336058 286008 336064
rect 285772 335368 285824 335374
rect 285772 335310 285824 335316
rect 285692 331186 285812 331214
rect 285588 331016 285640 331022
rect 285588 330958 285640 330964
rect 285404 326800 285456 326806
rect 285404 326742 285456 326748
rect 284944 326732 284996 326738
rect 284944 326674 284996 326680
rect 285784 316034 285812 331186
rect 286060 325174 286088 337742
rect 286336 335696 286364 338014
rect 286474 337770 286502 338028
rect 286244 335668 286364 335696
rect 286428 337742 286502 337770
rect 286566 337770 286594 338028
rect 286704 338014 286764 338042
rect 286566 337742 286640 337770
rect 286244 332314 286272 335668
rect 286324 335436 286376 335442
rect 286324 335378 286376 335384
rect 286232 332308 286284 332314
rect 286232 332250 286284 332256
rect 286048 325168 286100 325174
rect 286048 325110 286100 325116
rect 285692 316006 285812 316034
rect 284484 9104 284536 9110
rect 284484 9046 284536 9052
rect 284392 5500 284444 5506
rect 284392 5442 284444 5448
rect 285404 5092 285456 5098
rect 285404 5034 285456 5040
rect 285416 480 285444 5034
rect 285692 4214 285720 316006
rect 286336 5098 286364 335378
rect 286428 323678 286456 337742
rect 286612 337634 286640 337742
rect 286520 337606 286640 337634
rect 286520 335782 286548 337606
rect 286600 336524 286652 336530
rect 286600 336466 286652 336472
rect 286508 335776 286560 335782
rect 286508 335718 286560 335724
rect 286506 335472 286562 335481
rect 286506 335407 286562 335416
rect 286520 327962 286548 335407
rect 286612 334150 286640 336466
rect 286600 334144 286652 334150
rect 286600 334086 286652 334092
rect 286704 330954 286732 338014
rect 286842 337770 286870 338028
rect 286934 337872 286962 338028
rect 287072 338014 287132 338042
rect 286934 337844 287008 337872
rect 286796 337742 286870 337770
rect 286692 330948 286744 330954
rect 286692 330890 286744 330896
rect 286508 327956 286560 327962
rect 286508 327898 286560 327904
rect 286796 327826 286824 337742
rect 286980 336598 287008 337844
rect 286968 336592 287020 336598
rect 286968 336534 287020 336540
rect 286968 336048 287020 336054
rect 286968 335990 287020 335996
rect 286876 335368 286928 335374
rect 286876 335310 286928 335316
rect 286784 327820 286836 327826
rect 286784 327762 286836 327768
rect 286888 326602 286916 335310
rect 286980 334014 287008 335990
rect 286968 334008 287020 334014
rect 286968 333950 287020 333956
rect 287072 333606 287100 338014
rect 287210 337770 287238 338028
rect 287302 337906 287330 338028
rect 287440 338014 287500 338042
rect 287302 337878 287376 337906
rect 287210 337742 287284 337770
rect 287256 335578 287284 337742
rect 287348 336530 287376 337878
rect 287336 336524 287388 336530
rect 287336 336466 287388 336472
rect 287334 336016 287390 336025
rect 287334 335951 287390 335960
rect 287244 335572 287296 335578
rect 287244 335514 287296 335520
rect 287244 335436 287296 335442
rect 287244 335378 287296 335384
rect 287060 333600 287112 333606
rect 287060 333542 287112 333548
rect 287060 331900 287112 331906
rect 287060 331842 287112 331848
rect 286876 326596 286928 326602
rect 286876 326538 286928 326544
rect 286416 323672 286468 323678
rect 286416 323614 286468 323620
rect 287072 16574 287100 331842
rect 287256 323610 287284 335378
rect 287348 333810 287376 335951
rect 287336 333804 287388 333810
rect 287336 333746 287388 333752
rect 287440 332246 287468 338014
rect 287578 337770 287606 338028
rect 287670 337872 287698 338028
rect 287762 337940 287790 338028
rect 287900 338014 287960 338042
rect 287762 337912 287836 337940
rect 287670 337844 287744 337872
rect 287578 337742 287652 337770
rect 287520 335844 287572 335850
rect 287520 335786 287572 335792
rect 287532 334830 287560 335786
rect 287624 335510 287652 337742
rect 287716 336054 287744 337844
rect 287704 336048 287756 336054
rect 287704 335990 287756 335996
rect 287612 335504 287664 335510
rect 287612 335446 287664 335452
rect 287704 335368 287756 335374
rect 287704 335310 287756 335316
rect 287520 334824 287572 334830
rect 287520 334766 287572 334772
rect 287428 332240 287480 332246
rect 287428 332182 287480 332188
rect 287244 323604 287296 323610
rect 287244 323546 287296 323552
rect 287716 316034 287744 335310
rect 287808 330886 287836 337912
rect 287900 335442 287928 338014
rect 288038 337770 288066 338028
rect 288130 337872 288158 338028
rect 288268 338014 288328 338042
rect 288130 337844 288204 337872
rect 288038 337742 288112 337770
rect 288084 335850 288112 337742
rect 288072 335844 288124 335850
rect 288072 335786 288124 335792
rect 287980 335572 288032 335578
rect 287980 335514 288032 335520
rect 287888 335436 287940 335442
rect 287888 335378 287940 335384
rect 287992 331214 288020 335514
rect 288072 335504 288124 335510
rect 288072 335446 288124 335452
rect 288084 334506 288112 335446
rect 288176 335186 288204 337844
rect 288268 335374 288296 338014
rect 288406 337770 288434 338028
rect 288360 337742 288434 337770
rect 288498 337770 288526 338028
rect 288636 338014 288696 338042
rect 288498 337742 288572 337770
rect 288360 336025 288388 337742
rect 288346 336016 288402 336025
rect 288346 335951 288402 335960
rect 288256 335368 288308 335374
rect 288256 335310 288308 335316
rect 288176 335158 288296 335186
rect 288084 334478 288204 334506
rect 287992 331186 288112 331214
rect 287796 330880 287848 330886
rect 287796 330822 287848 330828
rect 288084 326534 288112 331186
rect 288072 326528 288124 326534
rect 288072 326470 288124 326476
rect 288176 325106 288204 334478
rect 288268 329458 288296 335158
rect 288544 332110 288572 337742
rect 288636 335510 288664 338014
rect 288774 337770 288802 338028
rect 288866 337872 288894 338028
rect 289004 338014 289064 338042
rect 288866 337844 288940 337872
rect 288774 337742 288848 337770
rect 288820 335714 288848 337742
rect 288808 335708 288860 335714
rect 288808 335650 288860 335656
rect 288912 335594 288940 337844
rect 288820 335566 288940 335594
rect 288624 335504 288676 335510
rect 288624 335446 288676 335452
rect 288820 333470 288848 335566
rect 289004 335442 289032 338014
rect 289142 337770 289170 338028
rect 289234 337872 289262 338028
rect 289372 338014 289432 338042
rect 289234 337844 289308 337872
rect 289142 337742 289216 337770
rect 289084 336456 289136 336462
rect 289084 336398 289136 336404
rect 288992 335436 289044 335442
rect 288992 335378 289044 335384
rect 288900 335368 288952 335374
rect 288900 335310 288952 335316
rect 288808 333464 288860 333470
rect 288808 333406 288860 333412
rect 288532 332104 288584 332110
rect 288532 332046 288584 332052
rect 288256 329452 288308 329458
rect 288256 329394 288308 329400
rect 288164 325100 288216 325106
rect 288164 325042 288216 325048
rect 288912 322250 288940 335310
rect 288992 326392 289044 326398
rect 288992 326334 289044 326340
rect 288900 322244 288952 322250
rect 288900 322186 288952 322192
rect 287624 316006 287744 316034
rect 287072 16546 287376 16574
rect 286324 5092 286376 5098
rect 286324 5034 286376 5040
rect 286600 5024 286652 5030
rect 286600 4966 286652 4972
rect 285680 4208 285732 4214
rect 285680 4150 285732 4156
rect 286612 480 286640 4966
rect 287348 490 287376 16546
rect 287624 13190 287652 316006
rect 287612 13184 287664 13190
rect 287612 13126 287664 13132
rect 289004 5506 289032 326334
rect 288992 5500 289044 5506
rect 288992 5442 289044 5448
rect 288992 4888 289044 4894
rect 288992 4830 289044 4836
rect 287624 598 287836 626
rect 287624 490 287652 598
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 462 287652 490
rect 287808 480 287836 598
rect 289004 480 289032 4830
rect 289096 4214 289124 336398
rect 289188 335646 289216 337742
rect 289176 335640 289228 335646
rect 289176 335582 289228 335588
rect 289280 330750 289308 337844
rect 289372 335374 289400 338014
rect 289510 337770 289538 338028
rect 289602 337906 289630 338028
rect 289740 338014 289800 338042
rect 289602 337878 289676 337906
rect 289510 337742 289584 337770
rect 289556 335986 289584 337742
rect 289544 335980 289596 335986
rect 289544 335922 289596 335928
rect 289452 335504 289504 335510
rect 289452 335446 289504 335452
rect 289360 335368 289412 335374
rect 289360 335310 289412 335316
rect 289268 330744 289320 330750
rect 289268 330686 289320 330692
rect 289464 326466 289492 335446
rect 289544 335436 289596 335442
rect 289544 335378 289596 335384
rect 289452 326460 289504 326466
rect 289452 326402 289504 326408
rect 289556 325038 289584 335378
rect 289648 329390 289676 337878
rect 289636 329384 289688 329390
rect 289636 329326 289688 329332
rect 289740 326398 289768 338014
rect 289878 337770 289906 338028
rect 289970 337906 289998 338028
rect 290108 338014 290168 338042
rect 289970 337878 290044 337906
rect 289878 337742 289952 337770
rect 289924 335510 289952 337742
rect 289912 335504 289964 335510
rect 289912 335446 289964 335452
rect 290016 334626 290044 337878
rect 290108 335374 290136 338014
rect 290246 337770 290274 338028
rect 290338 337906 290366 338028
rect 290338 337878 290412 337906
rect 290246 337742 290320 337770
rect 290292 336297 290320 337742
rect 290278 336288 290334 336297
rect 290278 336223 290334 336232
rect 290096 335368 290148 335374
rect 290096 335310 290148 335316
rect 290004 334620 290056 334626
rect 290004 334562 290056 334568
rect 290384 331974 290412 337878
rect 290522 337770 290550 338028
rect 290614 337958 290642 338028
rect 290602 337952 290654 337958
rect 290706 337940 290734 338028
rect 290844 338014 290904 338042
rect 290706 337912 290780 337940
rect 290602 337894 290654 337900
rect 290522 337742 290596 337770
rect 290372 331968 290424 331974
rect 290372 331910 290424 331916
rect 290568 326738 290596 337742
rect 290752 333402 290780 337912
rect 290740 333396 290792 333402
rect 290740 333338 290792 333344
rect 290556 326732 290608 326738
rect 290556 326674 290608 326680
rect 289728 326392 289780 326398
rect 289728 326334 289780 326340
rect 289544 325032 289596 325038
rect 289544 324974 289596 324980
rect 290844 324970 290872 338014
rect 290982 337770 291010 338028
rect 291074 337906 291102 338028
rect 291212 338014 291272 338042
rect 291074 337878 291148 337906
rect 290982 337742 291056 337770
rect 291028 335481 291056 337742
rect 291014 335472 291070 335481
rect 291014 335407 291070 335416
rect 290924 335368 290976 335374
rect 290924 335310 290976 335316
rect 290936 328030 290964 335310
rect 291120 330682 291148 337878
rect 291212 333334 291240 338014
rect 291350 337770 291378 338028
rect 291442 337929 291470 338028
rect 291534 337940 291562 338028
rect 291672 338014 291732 338042
rect 291428 337920 291484 337929
rect 291534 337912 291608 337940
rect 291428 337855 291484 337864
rect 291350 337742 291424 337770
rect 291396 336569 291424 337742
rect 291382 336560 291438 336569
rect 291382 336495 291438 336504
rect 291200 333328 291252 333334
rect 291200 333270 291252 333276
rect 291108 330676 291160 330682
rect 291108 330618 291160 330624
rect 291200 329112 291252 329118
rect 291200 329054 291252 329060
rect 290924 328024 290976 328030
rect 290924 327966 290976 327972
rect 290832 324964 290884 324970
rect 290832 324906 290884 324912
rect 291212 16574 291240 329054
rect 291580 323746 291608 337912
rect 291672 336161 291700 338014
rect 291810 337940 291838 338028
rect 291764 337912 291838 337940
rect 291902 337940 291930 338028
rect 292040 338014 292100 338042
rect 291902 337912 291976 337940
rect 291764 337770 291792 337912
rect 291764 337742 291884 337770
rect 291658 336152 291714 336161
rect 291658 336087 291714 336096
rect 291752 335368 291804 335374
rect 291752 335310 291804 335316
rect 291764 329186 291792 335310
rect 291856 329254 291884 337742
rect 291844 329248 291896 329254
rect 291844 329190 291896 329196
rect 291752 329180 291804 329186
rect 291752 329122 291804 329128
rect 291568 323740 291620 323746
rect 291568 323682 291620 323688
rect 291948 322318 291976 337912
rect 292040 334937 292068 338014
rect 292178 337906 292206 338028
rect 292132 337878 292206 337906
rect 292132 335374 292160 337878
rect 292270 337770 292298 338028
rect 292224 337742 292298 337770
rect 292408 338014 292468 338042
rect 292120 335368 292172 335374
rect 292120 335310 292172 335316
rect 292026 334928 292082 334937
rect 292026 334863 292082 334872
rect 292120 333736 292172 333742
rect 292120 333678 292172 333684
rect 292132 327758 292160 333678
rect 292120 327752 292172 327758
rect 292120 327694 292172 327700
rect 291936 322312 291988 322318
rect 291936 322254 291988 322260
rect 292224 321554 292252 337742
rect 292408 334801 292436 338014
rect 292546 337770 292574 338028
rect 292500 337742 292574 337770
rect 292638 337770 292666 338028
rect 292776 338014 292836 338042
rect 292638 337742 292712 337770
rect 292394 334792 292450 334801
rect 292394 334727 292450 334736
rect 292500 333742 292528 337742
rect 292684 335374 292712 337742
rect 292776 335714 292804 338014
rect 292914 337770 292942 338028
rect 293006 337906 293034 338028
rect 293144 338014 293204 338042
rect 293006 337878 293080 337906
rect 292914 337742 292988 337770
rect 292960 336938 292988 337742
rect 292948 336932 293000 336938
rect 292948 336874 293000 336880
rect 292764 335708 292816 335714
rect 292764 335650 292816 335656
rect 292580 335368 292632 335374
rect 292580 335310 292632 335316
rect 292672 335368 292724 335374
rect 292672 335310 292724 335316
rect 292592 333742 292620 335310
rect 292488 333736 292540 333742
rect 292488 333678 292540 333684
rect 292580 333736 292632 333742
rect 292580 333678 292632 333684
rect 292304 333328 292356 333334
rect 292304 333270 292356 333276
rect 292316 325242 292344 333270
rect 293052 331158 293080 337878
rect 293144 335617 293172 338014
rect 293282 337770 293310 338028
rect 293374 337906 293402 338028
rect 293374 337878 293448 337906
rect 293282 337742 293356 337770
rect 293130 335608 293186 335617
rect 293130 335543 293186 335552
rect 293040 331152 293092 331158
rect 293040 331094 293092 331100
rect 293328 330614 293356 337742
rect 293316 330608 293368 330614
rect 293316 330550 293368 330556
rect 292304 325236 292356 325242
rect 292304 325178 292356 325184
rect 293420 323814 293448 337878
rect 293558 337770 293586 338028
rect 293650 337890 293678 338028
rect 293742 337940 293770 338028
rect 293880 338014 293940 338042
rect 293742 337912 293816 337940
rect 293638 337884 293690 337890
rect 293638 337826 293690 337832
rect 293558 337742 293632 337770
rect 293604 335753 293632 337742
rect 293590 335744 293646 335753
rect 293590 335679 293646 335688
rect 293788 334676 293816 337912
rect 293880 335458 293908 338014
rect 294018 337770 294046 338028
rect 294110 337906 294138 338028
rect 294248 338014 294308 338042
rect 294110 337878 294184 337906
rect 294018 337742 294092 337770
rect 293880 335430 294000 335458
rect 293868 335368 293920 335374
rect 293868 335310 293920 335316
rect 293604 334648 293816 334676
rect 293604 326806 293632 334648
rect 293880 331214 293908 335310
rect 293972 334665 294000 335430
rect 293958 334656 294014 334665
rect 293958 334591 294014 334600
rect 293696 331186 293908 331214
rect 293696 328098 293724 331186
rect 294064 330546 294092 337742
rect 294156 336870 294184 337878
rect 294144 336864 294196 336870
rect 294144 336806 294196 336812
rect 294248 335442 294276 338014
rect 294386 337770 294414 338028
rect 294478 337958 294506 338028
rect 294466 337952 294518 337958
rect 294466 337894 294518 337900
rect 294662 337890 294690 338028
rect 294754 337906 294782 338028
rect 294860 338014 295104 338042
rect 294972 337952 295024 337958
rect 294650 337884 294702 337890
rect 294754 337878 294828 337906
rect 294972 337894 295024 337900
rect 294650 337826 294702 337832
rect 294386 337742 294736 337770
rect 294604 335912 294656 335918
rect 294604 335854 294656 335860
rect 294236 335436 294288 335442
rect 294236 335378 294288 335384
rect 294052 330540 294104 330546
rect 294052 330482 294104 330488
rect 293684 328092 293736 328098
rect 293684 328034 293736 328040
rect 293592 326800 293644 326806
rect 293592 326742 293644 326748
rect 293408 323808 293460 323814
rect 293408 323750 293460 323756
rect 292040 321526 292252 321554
rect 291212 16546 291424 16574
rect 289544 5500 289596 5506
rect 289544 5442 289596 5448
rect 289556 4894 289584 5442
rect 289544 4888 289596 4894
rect 289544 4830 289596 4836
rect 290188 4344 290240 4350
rect 290188 4286 290240 4292
rect 289084 4208 289136 4214
rect 289084 4150 289136 4156
rect 290200 480 290228 4286
rect 291396 480 291424 16546
rect 292040 13122 292068 321526
rect 292028 13116 292080 13122
rect 292028 13058 292080 13064
rect 294616 6798 294644 335854
rect 294708 8974 294736 337742
rect 294800 335374 294828 337878
rect 294880 337884 294932 337890
rect 294880 337826 294932 337832
rect 294892 335578 294920 337826
rect 294984 336802 295012 337894
rect 294972 336796 295024 336802
rect 294972 336738 295024 336744
rect 294972 336048 295024 336054
rect 294972 335990 295024 335996
rect 294880 335572 294932 335578
rect 294880 335514 294932 335520
rect 294880 335436 294932 335442
rect 294880 335378 294932 335384
rect 294788 335368 294840 335374
rect 294788 335310 294840 335316
rect 294788 330540 294840 330546
rect 294788 330482 294840 330488
rect 294800 9042 294828 330482
rect 294892 16574 294920 335378
rect 294984 20670 295012 335990
rect 294972 20664 295024 20670
rect 294972 20606 295024 20612
rect 294892 16546 295012 16574
rect 294788 9036 294840 9042
rect 294788 8978 294840 8984
rect 294696 8968 294748 8974
rect 294696 8910 294748 8916
rect 294604 6792 294656 6798
rect 294604 6734 294656 6740
rect 294984 4826 295012 16546
rect 292580 4820 292632 4826
rect 292580 4762 292632 4768
rect 294972 4820 295024 4826
rect 294972 4762 295024 4768
rect 292592 480 292620 4762
rect 293684 4276 293736 4282
rect 293684 4218 293736 4224
rect 293696 480 293724 4218
rect 294880 4208 294932 4214
rect 294880 4150 294932 4156
rect 294892 480 294920 4150
rect 295076 3369 295104 338014
rect 295168 335918 295196 340846
rect 295260 336054 295288 344986
rect 295522 337920 295578 337929
rect 295522 337855 295578 337864
rect 295248 336048 295300 336054
rect 295248 335990 295300 335996
rect 295156 335912 295208 335918
rect 295156 335854 295208 335860
rect 295248 335572 295300 335578
rect 295248 335514 295300 335520
rect 295156 335368 295208 335374
rect 295156 335310 295208 335316
rect 295168 3505 295196 335310
rect 295260 3641 295288 335514
rect 295432 335436 295484 335442
rect 295432 335378 295484 335384
rect 295340 334688 295392 334694
rect 295340 334630 295392 334636
rect 295246 3632 295302 3641
rect 295246 3567 295302 3576
rect 295154 3496 295210 3505
rect 295154 3431 295210 3440
rect 295062 3360 295118 3369
rect 295062 3295 295118 3304
rect 295352 626 295380 334630
rect 295444 4350 295472 335378
rect 295536 331906 295564 337855
rect 295708 335912 295760 335918
rect 295708 335854 295760 335860
rect 295524 331900 295576 331906
rect 295524 331842 295576 331848
rect 295720 316034 295748 335854
rect 295798 335608 295854 335617
rect 295798 335543 295854 335552
rect 295812 330614 295840 335543
rect 295800 330608 295852 330614
rect 295800 330550 295852 330556
rect 295536 316006 295748 316034
rect 295432 4344 295484 4350
rect 295432 4286 295484 4292
rect 295536 4282 295564 316006
rect 295996 206990 296024 379306
rect 302884 379160 302936 379166
rect 302884 379102 302936 379108
rect 300216 377868 300268 377874
rect 300216 377810 300268 377816
rect 298836 377800 298888 377806
rect 298836 377742 298888 377748
rect 298744 336728 298796 336734
rect 298744 336670 298796 336676
rect 296442 336560 296498 336569
rect 296442 336495 296498 336504
rect 296352 335368 296404 335374
rect 296352 335310 296404 335316
rect 296364 332178 296392 335310
rect 296456 333334 296484 336495
rect 296628 335776 296680 335782
rect 296628 335718 296680 335724
rect 298006 335744 298062 335753
rect 296536 335640 296588 335646
rect 296536 335582 296588 335588
rect 296548 334694 296576 335582
rect 296640 334830 296668 335718
rect 298006 335679 298062 335688
rect 296628 334824 296680 334830
rect 296628 334766 296680 334772
rect 296536 334688 296588 334694
rect 296536 334630 296588 334636
rect 296444 333328 296496 333334
rect 296444 333270 296496 333276
rect 298020 333266 298048 335679
rect 298192 335572 298244 335578
rect 298192 335514 298244 335520
rect 298204 333674 298232 335514
rect 298100 333668 298152 333674
rect 298100 333610 298152 333616
rect 298192 333668 298244 333674
rect 298192 333610 298244 333616
rect 298008 333260 298060 333266
rect 298008 333202 298060 333208
rect 296352 332172 296404 332178
rect 296352 332114 296404 332120
rect 295984 206984 296036 206990
rect 295984 206926 296036 206932
rect 297272 9376 297324 9382
rect 297272 9318 297324 9324
rect 295524 4276 295576 4282
rect 295524 4218 295576 4224
rect 295352 598 295656 626
rect 295628 490 295656 598
rect 295904 598 296116 626
rect 295904 490 295932 598
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 295628 462 295932 490
rect 296088 480 296116 598
rect 297284 480 297312 9318
rect 298112 490 298140 333610
rect 298756 5030 298784 336670
rect 298848 245614 298876 377742
rect 299938 336288 299994 336297
rect 299938 336223 299994 336232
rect 299480 335844 299532 335850
rect 299480 335786 299532 335792
rect 299492 334762 299520 335786
rect 299388 334756 299440 334762
rect 299388 334698 299440 334704
rect 299480 334756 299532 334762
rect 299480 334698 299532 334704
rect 299400 334642 299428 334698
rect 299400 334614 299520 334642
rect 298836 245608 298888 245614
rect 298836 245550 298888 245556
rect 299492 16574 299520 334614
rect 299952 330818 299980 336223
rect 300124 333532 300176 333538
rect 300124 333474 300176 333480
rect 299940 330812 299992 330818
rect 299940 330754 299992 330760
rect 299492 16546 299704 16574
rect 298744 5024 298796 5030
rect 298744 4966 298796 4972
rect 298296 598 298508 626
rect 298296 490 298324 598
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 462 298324 490
rect 298480 480 298508 598
rect 299676 480 299704 16546
rect 300136 2854 300164 333474
rect 300228 299470 300256 377810
rect 302896 353258 302924 379102
rect 304264 379024 304316 379030
rect 304264 378966 304316 378972
rect 302884 353252 302936 353258
rect 302884 353194 302936 353200
rect 303252 335980 303304 335986
rect 303252 335922 303304 335928
rect 302240 334008 302292 334014
rect 302240 333950 302292 333956
rect 300216 299464 300268 299470
rect 300216 299406 300268 299412
rect 302252 16574 302280 333950
rect 303264 333538 303292 335922
rect 304172 335844 304224 335850
rect 304172 335786 304224 335792
rect 303252 333532 303304 333538
rect 303252 333474 303304 333480
rect 304184 329322 304212 335786
rect 304172 329316 304224 329322
rect 304172 329258 304224 329264
rect 304276 193186 304304 378966
rect 307116 378888 307168 378894
rect 307116 378830 307168 378836
rect 305644 377664 305696 377670
rect 305644 377606 305696 377612
rect 305000 331424 305052 331430
rect 305000 331366 305052 331372
rect 304264 193180 304316 193186
rect 304264 193122 304316 193128
rect 305012 16574 305040 331366
rect 305656 233238 305684 377606
rect 306380 334076 306432 334082
rect 306380 334018 306432 334024
rect 305644 233232 305696 233238
rect 305644 233174 305696 233180
rect 302252 16546 303200 16574
rect 305012 16546 305592 16574
rect 300768 9308 300820 9314
rect 300768 9250 300820 9256
rect 300124 2848 300176 2854
rect 300124 2790 300176 2796
rect 300780 480 300808 9250
rect 301964 2848 302016 2854
rect 301964 2790 302016 2796
rect 301976 480 302004 2790
rect 303172 480 303200 16546
rect 304356 9240 304408 9246
rect 304356 9182 304408 9188
rect 304368 480 304396 9182
rect 305564 480 305592 16546
rect 306392 490 306420 334018
rect 307024 332716 307076 332722
rect 307024 332658 307076 332664
rect 307036 2854 307064 332658
rect 307128 273222 307156 378830
rect 314016 378820 314068 378826
rect 314016 378762 314068 378768
rect 309784 377596 309836 377602
rect 309784 377538 309836 377544
rect 309140 334144 309192 334150
rect 309140 334086 309192 334092
rect 307116 273216 307168 273222
rect 307116 273158 307168 273164
rect 309152 16574 309180 334086
rect 309796 325650 309824 377538
rect 313280 334212 313332 334218
rect 313280 334154 313332 334160
rect 310520 332784 310572 332790
rect 310520 332726 310572 332732
rect 309784 325644 309836 325650
rect 309784 325586 309836 325592
rect 310532 16574 310560 332726
rect 311900 325440 311952 325446
rect 311900 325382 311952 325388
rect 311912 16574 311940 325382
rect 313292 16574 313320 334154
rect 313924 331492 313976 331498
rect 313924 331434 313976 331440
rect 309152 16546 309824 16574
rect 310532 16546 311480 16574
rect 311912 16546 312216 16574
rect 313292 16546 313872 16574
rect 309048 5092 309100 5098
rect 309048 5034 309100 5040
rect 307024 2848 307076 2854
rect 307024 2790 307076 2796
rect 307944 2848 307996 2854
rect 307944 2790 307996 2796
rect 306576 598 306788 626
rect 306576 490 306604 598
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306392 462 306604 490
rect 306760 480 306788 598
rect 307956 480 307984 2790
rect 309060 480 309088 5034
rect 309796 490 309824 16546
rect 310072 598 310284 626
rect 310072 490 310100 598
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 462 310100 490
rect 310256 480 310284 598
rect 311452 480 311480 16546
rect 312188 490 312216 16546
rect 312464 598 312676 626
rect 312464 490 312492 598
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 462 312492 490
rect 312648 480 312676 598
rect 313844 480 313872 16546
rect 313936 2854 313964 331434
rect 314028 259418 314056 378762
rect 318064 378752 318116 378758
rect 318064 378694 318116 378700
rect 316684 377256 316736 377262
rect 316684 377198 316736 377204
rect 316040 334280 316092 334286
rect 316040 334222 316092 334228
rect 314016 259412 314068 259418
rect 314016 259354 314068 259360
rect 316052 2854 316080 334222
rect 316696 313274 316724 377198
rect 318076 365702 318104 378694
rect 580172 378480 580224 378486
rect 580170 378448 580172 378457
rect 580224 378448 580226 378457
rect 580170 378383 580226 378392
rect 318064 365696 318116 365702
rect 318064 365638 318116 365644
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 349160 337680 349212 337686
rect 349160 337622 349212 337628
rect 320824 336660 320876 336666
rect 320824 336602 320876 336608
rect 317420 330268 317472 330274
rect 317420 330210 317472 330216
rect 316684 313268 316736 313274
rect 316684 313210 316736 313216
rect 317432 16574 317460 330210
rect 317432 16546 318104 16574
rect 316224 15904 316276 15910
rect 316224 15846 316276 15852
rect 313924 2848 313976 2854
rect 313924 2790 313976 2796
rect 315028 2848 315080 2854
rect 315028 2790 315080 2796
rect 316040 2848 316092 2854
rect 316040 2790 316092 2796
rect 315040 480 315068 2790
rect 316236 480 316264 15846
rect 317328 2848 317380 2854
rect 317328 2790 317380 2796
rect 317340 480 317368 2790
rect 318076 490 318104 16546
rect 320836 5030 320864 336602
rect 322204 336592 322256 336598
rect 322204 336534 322256 336540
rect 321560 332852 321612 332858
rect 321560 332794 321612 332800
rect 321572 16574 321600 332794
rect 321572 16546 322152 16574
rect 320824 5024 320876 5030
rect 320824 4966 320876 4972
rect 319720 4956 319772 4962
rect 319720 4898 319772 4904
rect 320916 4956 320968 4962
rect 320916 4898 320968 4904
rect 318352 598 318564 626
rect 318352 490 318380 598
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 462 318380 490
rect 318536 480 318564 598
rect 319732 480 319760 4898
rect 320928 480 320956 4898
rect 322124 480 322152 16546
rect 322216 4962 322244 336534
rect 323676 336524 323728 336530
rect 323676 336466 323728 336472
rect 323584 336388 323636 336394
rect 323584 336330 323636 336336
rect 322940 325372 322992 325378
rect 322940 325314 322992 325320
rect 322204 4956 322256 4962
rect 322204 4898 322256 4904
rect 322952 490 322980 325314
rect 323596 15570 323624 336330
rect 323688 289134 323716 336466
rect 331864 336456 331916 336462
rect 331864 336398 331916 336404
rect 327722 336152 327778 336161
rect 327722 336087 327778 336096
rect 324962 336016 325018 336025
rect 324962 335951 325018 335960
rect 324320 334348 324372 334354
rect 324320 334290 324372 334296
rect 323676 289128 323728 289134
rect 323676 289070 323728 289076
rect 323584 15564 323636 15570
rect 323584 15506 323636 15512
rect 324332 6914 324360 334290
rect 324412 331560 324464 331566
rect 324412 331502 324464 331508
rect 324424 11694 324452 331502
rect 324976 177342 325004 335951
rect 324964 177336 325016 177342
rect 324964 177278 325016 177284
rect 327736 17270 327764 336087
rect 328460 330336 328512 330342
rect 328460 330278 328512 330284
rect 327724 17264 327776 17270
rect 327724 17206 327776 17212
rect 328472 16574 328500 330278
rect 329840 323944 329892 323950
rect 329840 323886 329892 323892
rect 329852 16574 329880 323886
rect 328472 16546 328776 16574
rect 329852 16546 330432 16574
rect 328000 15564 328052 15570
rect 328000 15506 328052 15512
rect 324412 11688 324464 11694
rect 324412 11630 324464 11636
rect 325608 11688 325660 11694
rect 325608 11630 325660 11636
rect 324332 6886 324452 6914
rect 323136 598 323348 626
rect 323136 490 323164 598
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 322952 462 323164 490
rect 323320 480 323348 598
rect 324424 480 324452 6886
rect 325620 480 325648 11630
rect 326804 9172 326856 9178
rect 326804 9114 326856 9120
rect 326816 480 326844 9114
rect 328012 480 328040 15506
rect 328748 490 328776 16546
rect 329024 598 329236 626
rect 329024 490 329052 598
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 328748 462 329052 490
rect 329208 480 329236 598
rect 330404 480 330432 16546
rect 331588 5704 331640 5710
rect 331588 5646 331640 5652
rect 331600 480 331628 5646
rect 331876 5098 331904 336398
rect 336004 336320 336056 336326
rect 336004 336262 336056 336268
rect 333980 334416 334032 334422
rect 333980 334358 334032 334364
rect 331956 332920 332008 332926
rect 331956 332862 332008 332868
rect 331864 5092 331916 5098
rect 331864 5034 331916 5040
rect 331968 2854 331996 332862
rect 333992 2854 334020 334358
rect 335360 331628 335412 331634
rect 335360 331570 335412 331576
rect 335372 16574 335400 331570
rect 335372 16546 335952 16574
rect 335084 5772 335136 5778
rect 335084 5714 335136 5720
rect 331956 2848 332008 2854
rect 331956 2790 332008 2796
rect 332692 2848 332744 2854
rect 332692 2790 332744 2796
rect 333980 2848 334032 2854
rect 333980 2790 334032 2796
rect 332704 480 332732 2790
rect 333888 2780 333940 2786
rect 333888 2722 333940 2728
rect 333900 480 333928 2722
rect 335096 480 335124 5714
rect 335924 3482 335952 16546
rect 336016 5166 336044 336262
rect 338120 331696 338172 331702
rect 338120 331638 338172 331644
rect 336004 5160 336056 5166
rect 336004 5102 336056 5108
rect 335924 3454 336320 3482
rect 336292 480 336320 3454
rect 338132 2854 338160 331638
rect 342904 330404 342956 330410
rect 342904 330346 342956 330352
rect 340880 328976 340932 328982
rect 340880 328918 340932 328924
rect 340892 16574 340920 328918
rect 342916 16574 342944 330346
rect 340892 16546 341012 16574
rect 342916 16546 343036 16574
rect 339500 9784 339552 9790
rect 339500 9726 339552 9732
rect 338672 5840 338724 5846
rect 338672 5782 338724 5788
rect 337476 2848 337528 2854
rect 337476 2790 337528 2796
rect 338120 2848 338172 2854
rect 338120 2790 338172 2796
rect 337488 480 337516 2790
rect 338684 480 338712 5782
rect 339512 490 339540 9726
rect 339696 598 339908 626
rect 339696 490 339724 598
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339512 462 339724 490
rect 339880 480 339908 598
rect 340984 480 341012 16546
rect 342904 9852 342956 9858
rect 342904 9794 342956 9800
rect 342168 5908 342220 5914
rect 342168 5850 342220 5856
rect 342180 480 342208 5850
rect 342916 490 342944 9794
rect 343008 2854 343036 16546
rect 346952 9920 347004 9926
rect 346952 9862 347004 9868
rect 345756 5976 345808 5982
rect 345756 5918 345808 5924
rect 342996 2848 343048 2854
rect 342996 2790 343048 2796
rect 344560 2848 344612 2854
rect 344560 2790 344612 2796
rect 343192 598 343404 626
rect 343192 490 343220 598
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 462 343220 490
rect 343376 480 343404 598
rect 344572 480 344600 2790
rect 345768 480 345796 5918
rect 346964 480 346992 9862
rect 349172 2854 349200 337622
rect 360844 337612 360896 337618
rect 360844 337554 360896 337560
rect 351920 334484 351972 334490
rect 351920 334426 351972 334432
rect 350448 9988 350500 9994
rect 350448 9930 350500 9936
rect 349252 6044 349304 6050
rect 349252 5986 349304 5992
rect 348056 2848 348108 2854
rect 348056 2790 348108 2796
rect 349160 2848 349212 2854
rect 349160 2790 349212 2796
rect 348068 480 348096 2790
rect 349264 480 349292 5986
rect 350460 480 350488 9930
rect 351932 3482 351960 334426
rect 353944 332988 353996 332994
rect 353944 332930 353996 332936
rect 353576 10056 353628 10062
rect 353576 9998 353628 10004
rect 352840 6112 352892 6118
rect 352840 6054 352892 6060
rect 351656 3454 351960 3482
rect 351656 480 351684 3454
rect 352852 480 352880 6054
rect 353588 490 353616 9998
rect 353956 2854 353984 332930
rect 357440 331764 357492 331770
rect 357440 331706 357492 331712
rect 356336 6724 356388 6730
rect 356336 6666 356388 6672
rect 353944 2848 353996 2854
rect 353944 2790 353996 2796
rect 355232 2848 355284 2854
rect 355232 2790 355284 2796
rect 353864 598 354076 626
rect 353864 490 353892 598
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 353588 462 353892 490
rect 354048 480 354076 598
rect 355244 480 355272 2790
rect 356348 480 356376 6666
rect 357452 2854 357480 331706
rect 360752 10192 360804 10198
rect 360752 10134 360804 10140
rect 357532 10124 357584 10130
rect 357532 10066 357584 10072
rect 357440 2848 357492 2854
rect 357440 2790 357492 2796
rect 357544 480 357572 10066
rect 359924 6656 359976 6662
rect 359924 6598 359976 6604
rect 358728 2848 358780 2854
rect 358728 2790 358780 2796
rect 358740 480 358768 2790
rect 359936 480 359964 6598
rect 360764 1986 360792 10134
rect 360856 2854 360884 337554
rect 367100 337544 367152 337550
rect 367100 337486 367152 337492
rect 364616 10260 364668 10266
rect 364616 10202 364668 10208
rect 363512 6588 363564 6594
rect 363512 6530 363564 6536
rect 360844 2848 360896 2854
rect 360844 2790 360896 2796
rect 362316 2848 362368 2854
rect 362316 2790 362368 2796
rect 360764 1958 361160 1986
rect 361132 480 361160 1958
rect 362328 480 362356 2790
rect 363524 480 363552 6530
rect 364628 480 364656 10202
rect 367008 6520 367060 6526
rect 367008 6462 367060 6468
rect 365812 2848 365864 2854
rect 365812 2790 365864 2796
rect 365824 480 365852 2790
rect 367020 480 367048 6462
rect 367112 2854 367140 337486
rect 369860 337476 369912 337482
rect 369860 337418 369912 337424
rect 367744 11008 367796 11014
rect 367744 10950 367796 10956
rect 367100 2848 367152 2854
rect 367100 2790 367152 2796
rect 367756 490 367784 10950
rect 369872 2854 369900 337418
rect 425704 337408 425756 337414
rect 425704 337350 425756 337356
rect 376024 336252 376076 336258
rect 376024 336194 376076 336200
rect 371884 334552 371936 334558
rect 371884 334494 371936 334500
rect 371240 10940 371292 10946
rect 371240 10882 371292 10888
rect 370596 6452 370648 6458
rect 370596 6394 370648 6400
rect 369400 2848 369452 2854
rect 369400 2790 369452 2796
rect 369860 2848 369912 2854
rect 369860 2790 369912 2796
rect 368032 598 368244 626
rect 368032 490 368060 598
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 462 368060 490
rect 368216 480 368244 598
rect 369412 480 369440 2790
rect 370608 480 370636 6394
rect 371252 490 371280 10882
rect 371896 2854 371924 334494
rect 375380 330472 375432 330478
rect 375380 330414 375432 330420
rect 374000 10872 374052 10878
rect 374000 10814 374052 10820
rect 374012 2854 374040 10814
rect 375392 6914 375420 330414
rect 376036 16574 376064 336194
rect 393964 336184 394016 336190
rect 393964 336126 394016 336132
rect 387800 335300 387852 335306
rect 387800 335242 387852 335248
rect 385684 331832 385736 331838
rect 385684 331774 385736 331780
rect 378784 329044 378836 329050
rect 378784 328986 378836 328992
rect 376036 16546 376156 16574
rect 375392 6886 376064 6914
rect 374092 6384 374144 6390
rect 374092 6326 374144 6332
rect 371884 2848 371936 2854
rect 371884 2790 371936 2796
rect 372896 2848 372948 2854
rect 372896 2790 372948 2796
rect 374000 2848 374052 2854
rect 374000 2790 374052 2796
rect 371528 598 371740 626
rect 371528 490 371556 598
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371252 462 371556 490
rect 371712 480 371740 598
rect 372908 480 372936 2790
rect 374104 480 374132 6326
rect 375288 2848 375340 2854
rect 375288 2790 375340 2796
rect 375300 480 375328 2790
rect 376036 490 376064 6886
rect 376128 5234 376156 16546
rect 378416 10804 378468 10810
rect 378416 10746 378468 10752
rect 377680 6316 377732 6322
rect 377680 6258 377732 6264
rect 376116 5228 376168 5234
rect 376116 5170 376168 5176
rect 376312 598 376524 626
rect 376312 490 376340 598
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 462 376340 490
rect 376496 480 376524 598
rect 377692 480 377720 6258
rect 378428 490 378456 10746
rect 378796 2854 378824 328986
rect 382280 328432 382332 328438
rect 382280 328374 382332 328380
rect 381176 6248 381228 6254
rect 381176 6190 381228 6196
rect 378784 2848 378836 2854
rect 378784 2790 378836 2796
rect 379980 2848 380032 2854
rect 379980 2790 380032 2796
rect 378704 598 378916 626
rect 378704 490 378732 598
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378428 462 378732 490
rect 378888 480 378916 598
rect 379992 480 380020 2790
rect 381188 480 381216 6190
rect 382292 2854 382320 328374
rect 382372 10736 382424 10742
rect 382372 10678 382424 10684
rect 382280 2848 382332 2854
rect 382280 2790 382332 2796
rect 382384 480 382412 10678
rect 385592 10668 385644 10674
rect 385592 10610 385644 10616
rect 384764 6180 384816 6186
rect 384764 6122 384816 6128
rect 383568 2848 383620 2854
rect 383568 2790 383620 2796
rect 383580 480 383608 2790
rect 384776 480 384804 6122
rect 385604 2666 385632 10610
rect 385696 2854 385724 331774
rect 385684 2848 385736 2854
rect 385684 2790 385736 2796
rect 387156 2848 387208 2854
rect 387156 2790 387208 2796
rect 385604 2638 386000 2666
rect 385972 480 386000 2638
rect 387168 480 387196 2790
rect 387812 490 387840 335242
rect 389824 329792 389876 329798
rect 389824 329734 389876 329740
rect 389456 10600 389508 10606
rect 389456 10542 389508 10548
rect 388088 598 388300 626
rect 388088 490 388116 598
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 387812 462 388116 490
rect 388272 480 388300 598
rect 389468 480 389496 10542
rect 389836 2854 389864 329734
rect 392584 328364 392636 328370
rect 392584 328306 392636 328312
rect 392596 16574 392624 328306
rect 392596 16546 392716 16574
rect 392584 10532 392636 10538
rect 392584 10474 392636 10480
rect 391848 5160 391900 5166
rect 391848 5102 391900 5108
rect 389824 2848 389876 2854
rect 389824 2790 389876 2796
rect 390652 2848 390704 2854
rect 390652 2790 390704 2796
rect 390664 480 390692 2790
rect 391860 480 391888 5102
rect 392596 490 392624 10474
rect 392688 2854 392716 16546
rect 393976 5166 394004 336126
rect 394700 335232 394752 335238
rect 394700 335174 394752 335180
rect 394712 16574 394740 335174
rect 414664 335164 414716 335170
rect 414664 335106 414716 335112
rect 405740 333192 405792 333198
rect 405740 333134 405792 333140
rect 398840 333056 398892 333062
rect 398840 332998 398892 333004
rect 396724 326936 396776 326942
rect 396724 326878 396776 326884
rect 394712 16546 395384 16574
rect 393964 5160 394016 5166
rect 393964 5102 394016 5108
rect 392676 2848 392728 2854
rect 392676 2790 392728 2796
rect 394240 2848 394292 2854
rect 394240 2790 394292 2796
rect 392872 598 393084 626
rect 392872 490 392900 598
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 462 392900 490
rect 393056 480 393084 598
rect 394252 480 394280 2790
rect 395356 480 395384 16546
rect 396080 10464 396132 10470
rect 396080 10406 396132 10412
rect 396092 490 396120 10406
rect 396736 2922 396764 326878
rect 398852 16574 398880 332998
rect 400220 325304 400272 325310
rect 400220 325246 400272 325252
rect 400232 16574 400260 325246
rect 403624 323876 403676 323882
rect 403624 323818 403676 323824
rect 398852 16546 398972 16574
rect 400232 16546 400904 16574
rect 396724 2916 396776 2922
rect 396724 2858 396776 2864
rect 397736 2916 397788 2922
rect 397736 2858 397788 2864
rect 396368 598 396580 626
rect 396368 490 396396 598
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 462 396396 490
rect 396552 480 396580 598
rect 397748 480 397776 2858
rect 398944 480 398972 16546
rect 400128 10396 400180 10402
rect 400128 10338 400180 10344
rect 400140 480 400168 10338
rect 400876 490 400904 16546
rect 403532 10328 403584 10334
rect 403532 10270 403584 10276
rect 402520 5228 402572 5234
rect 402520 5170 402572 5176
rect 401152 598 401364 626
rect 401152 490 401180 598
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 462 401180 490
rect 401336 480 401364 598
rect 402532 480 402560 5170
rect 403544 2802 403572 10270
rect 403636 2922 403664 323818
rect 405752 16574 405780 333134
rect 412640 333124 412692 333130
rect 412640 333066 412692 333072
rect 407120 329724 407172 329730
rect 407120 329666 407172 329672
rect 405752 16546 406056 16574
rect 403624 2916 403676 2922
rect 403624 2858 403676 2864
rect 404820 2916 404872 2922
rect 404820 2858 404872 2864
rect 403544 2774 403664 2802
rect 403636 480 403664 2774
rect 404832 480 404860 2858
rect 406028 480 406056 16546
rect 407132 6914 407160 329666
rect 409880 329656 409932 329662
rect 409880 329598 409932 329604
rect 407212 322380 407264 322386
rect 407212 322322 407264 322328
rect 407224 11694 407252 322322
rect 409892 16574 409920 329598
rect 409892 16546 410840 16574
rect 407212 11688 407264 11694
rect 407212 11630 407264 11636
rect 408408 11688 408460 11694
rect 408408 11630 408460 11636
rect 407132 6886 407252 6914
rect 407224 480 407252 6886
rect 408420 480 408448 11630
rect 409604 5160 409656 5166
rect 409604 5102 409656 5108
rect 409616 480 409644 5102
rect 410812 480 410840 16546
rect 411904 2848 411956 2854
rect 411904 2790 411956 2796
rect 411916 480 411944 2790
rect 412652 490 412680 333066
rect 414020 328296 414072 328302
rect 414020 328238 414072 328244
rect 414032 16574 414060 328238
rect 414032 16546 414336 16574
rect 412928 598 413140 626
rect 412928 490 412956 598
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 462 412956 490
rect 413112 480 413140 598
rect 414308 480 414336 16546
rect 414676 3194 414704 335106
rect 418804 333940 418856 333946
rect 418804 333882 418856 333888
rect 416780 328228 416832 328234
rect 416780 328170 416832 328176
rect 416792 16574 416820 328170
rect 416792 16546 417464 16574
rect 414664 3188 414716 3194
rect 414664 3130 414716 3136
rect 416688 3188 416740 3194
rect 416688 3130 416740 3136
rect 415492 3052 415544 3058
rect 415492 2994 415544 3000
rect 415504 480 415532 2994
rect 416700 480 416728 3130
rect 417436 490 417464 16546
rect 418816 3126 418844 333882
rect 423680 333872 423732 333878
rect 423680 333814 423732 333820
rect 420920 328160 420972 328166
rect 420920 328102 420972 328108
rect 418804 3120 418856 3126
rect 418804 3062 418856 3068
rect 420184 3120 420236 3126
rect 420184 3062 420236 3068
rect 418988 2848 419040 2854
rect 418988 2790 419040 2796
rect 417712 598 417924 626
rect 417712 490 417740 598
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 462 417740 490
rect 417896 480 417924 598
rect 419000 480 419028 2790
rect 420196 480 420224 3062
rect 420932 490 420960 328102
rect 423692 6914 423720 333814
rect 423772 326868 423824 326874
rect 423772 326810 423824 326816
rect 423784 11694 423812 326810
rect 423772 11688 423824 11694
rect 423772 11630 423824 11636
rect 424968 11688 425020 11694
rect 424968 11630 425020 11636
rect 423692 6886 423812 6914
rect 422576 2984 422628 2990
rect 422576 2926 422628 2932
rect 421208 598 421420 626
rect 421208 490 421236 598
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 420932 462 421236 490
rect 421392 480 421420 598
rect 422588 480 422616 2926
rect 423784 480 423812 6886
rect 424980 480 425008 11630
rect 425716 3330 425744 337350
rect 427820 337340 427872 337346
rect 427820 337282 427872 337288
rect 427832 16574 427860 337282
rect 432052 337272 432104 337278
rect 432052 337214 432104 337220
rect 430580 332580 430632 332586
rect 430580 332522 430632 332528
rect 430592 16574 430620 332522
rect 427832 16546 428504 16574
rect 430592 16546 430896 16574
rect 425704 3324 425756 3330
rect 425704 3266 425756 3272
rect 427268 3324 427320 3330
rect 427268 3266 427320 3272
rect 426164 3052 426216 3058
rect 426164 2994 426216 3000
rect 426176 480 426204 2994
rect 427280 480 427308 3266
rect 428476 480 428504 16546
rect 429660 3120 429712 3126
rect 429660 3062 429712 3068
rect 429672 480 429700 3062
rect 430868 480 430896 16546
rect 432064 480 432092 337214
rect 436744 337204 436796 337210
rect 436744 337146 436796 337152
rect 432604 335096 432656 335102
rect 432604 335038 432656 335044
rect 432616 3398 432644 335038
rect 434720 331220 434772 331226
rect 434720 331162 434772 331168
rect 434732 16574 434760 331162
rect 434732 16546 435128 16574
rect 432604 3392 432656 3398
rect 432604 3334 432656 3340
rect 434444 3392 434496 3398
rect 434444 3334 434496 3340
rect 433248 3256 433300 3262
rect 433248 3198 433300 3204
rect 433260 480 433288 3198
rect 434456 480 434484 3334
rect 435100 490 435128 16546
rect 436756 3398 436784 337146
rect 468484 337136 468536 337142
rect 468484 337078 468536 337084
rect 465172 333804 465224 333810
rect 465172 333746 465224 333752
rect 450544 331152 450596 331158
rect 450544 331094 450596 331100
rect 438860 329588 438912 329594
rect 438860 329530 438912 329536
rect 438872 16574 438900 329530
rect 443644 326800 443696 326806
rect 443644 326742 443696 326748
rect 438872 16546 439176 16574
rect 436744 3392 436796 3398
rect 436744 3334 436796 3340
rect 437940 3392 437992 3398
rect 437940 3334 437992 3340
rect 436744 3256 436796 3262
rect 436744 3198 436796 3204
rect 435376 598 435588 626
rect 435376 490 435404 598
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435100 462 435404 490
rect 435560 480 435588 598
rect 436756 480 436784 3198
rect 437952 480 437980 3334
rect 439148 480 439176 16546
rect 442632 12164 442684 12170
rect 442632 12106 442684 12112
rect 441528 8016 441580 8022
rect 441528 7958 441580 7964
rect 440332 4140 440384 4146
rect 440332 4082 440384 4088
rect 440344 480 440372 4082
rect 441540 480 441568 7958
rect 442644 480 442672 12106
rect 443656 4078 443684 326742
rect 447784 323808 447836 323814
rect 447784 323750 447836 323756
rect 445760 12096 445812 12102
rect 445760 12038 445812 12044
rect 445024 7948 445076 7954
rect 445024 7890 445076 7896
rect 443644 4072 443696 4078
rect 443644 4014 443696 4020
rect 443828 3324 443880 3330
rect 443828 3266 443880 3272
rect 443840 480 443868 3266
rect 445036 480 445064 7890
rect 445772 490 445800 12038
rect 447416 4004 447468 4010
rect 447416 3946 447468 3952
rect 446048 598 446260 626
rect 446048 490 446076 598
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 462 446076 490
rect 446232 480 446260 598
rect 447428 480 447456 3946
rect 447796 3942 447824 323750
rect 448520 12028 448572 12034
rect 448520 11970 448572 11976
rect 447784 3936 447836 3942
rect 447784 3878 447836 3884
rect 448532 3398 448560 11970
rect 448612 7880 448664 7886
rect 448612 7822 448664 7828
rect 448520 3392 448572 3398
rect 448520 3334 448572 3340
rect 448624 480 448652 7822
rect 450556 4010 450584 331094
rect 453304 328092 453356 328098
rect 453304 328034 453356 328040
rect 453212 11960 453264 11966
rect 453212 11902 453264 11908
rect 452108 7812 452160 7818
rect 452108 7754 452160 7760
rect 450084 4004 450136 4010
rect 450084 3946 450136 3952
rect 450544 4004 450596 4010
rect 450544 3946 450596 3952
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 449820 480 449848 3334
rect 450096 2854 450124 3946
rect 450084 2848 450136 2854
rect 450084 2790 450136 2796
rect 450912 2848 450964 2854
rect 450912 2790 450964 2796
rect 450924 480 450952 2790
rect 452120 480 452148 7754
rect 453224 3482 453252 11902
rect 453316 4146 453344 328034
rect 464344 328024 464396 328030
rect 464344 327966 464396 327972
rect 461584 326732 461636 326738
rect 461584 326674 461636 326680
rect 457444 325236 457496 325242
rect 457444 325178 457496 325184
rect 454684 323740 454736 323746
rect 454684 323682 454736 323688
rect 453304 4140 453356 4146
rect 453304 4082 453356 4088
rect 454696 3806 454724 323682
rect 456892 11892 456944 11898
rect 456892 11834 456944 11840
rect 455696 7744 455748 7750
rect 455696 7686 455748 7692
rect 454500 3800 454552 3806
rect 454500 3742 454552 3748
rect 454684 3800 454736 3806
rect 454684 3742 454736 3748
rect 453224 3454 453344 3482
rect 453316 480 453344 3454
rect 454512 480 454540 3742
rect 455708 480 455736 7686
rect 456904 480 456932 11834
rect 457456 3806 457484 325178
rect 461596 16574 461624 326674
rect 461596 16546 461716 16574
rect 459928 11824 459980 11830
rect 459928 11766 459980 11772
rect 459192 7676 459244 7682
rect 459192 7618 459244 7624
rect 457444 3800 457496 3806
rect 457444 3742 457496 3748
rect 458088 3392 458140 3398
rect 458088 3334 458140 3340
rect 458100 480 458128 3334
rect 459204 480 459232 7618
rect 459940 490 459968 11766
rect 461688 3738 461716 16546
rect 463976 11756 464028 11762
rect 463976 11698 464028 11704
rect 462780 7608 462832 7614
rect 462780 7550 462832 7556
rect 461584 3732 461636 3738
rect 461584 3674 461636 3680
rect 461676 3732 461728 3738
rect 461676 3674 461728 3680
rect 460216 598 460428 626
rect 460216 490 460244 598
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 462 460244 490
rect 460400 480 460428 598
rect 461596 480 461624 3674
rect 462792 480 462820 7550
rect 463988 480 464016 11698
rect 464356 3398 464384 327966
rect 465184 16574 465212 333746
rect 466460 327956 466512 327962
rect 466460 327898 466512 327904
rect 466472 16574 466500 327898
rect 465184 16546 465856 16574
rect 466472 16546 467512 16574
rect 465172 3664 465224 3670
rect 465172 3606 465224 3612
rect 464344 3392 464396 3398
rect 464344 3334 464396 3340
rect 465184 480 465212 3606
rect 465828 490 465856 16546
rect 466104 598 466316 626
rect 466104 490 466132 598
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 462 466132 490
rect 466288 480 466316 598
rect 467484 480 467512 16546
rect 468496 3602 468524 337078
rect 470600 337068 470652 337074
rect 470600 337010 470652 337016
rect 468668 3664 468720 3670
rect 468668 3606 468720 3612
rect 468484 3596 468536 3602
rect 468484 3538 468536 3544
rect 468680 480 468708 3606
rect 469864 3596 469916 3602
rect 469864 3538 469916 3544
rect 469876 480 469904 3538
rect 470612 490 470640 337010
rect 472624 337000 472676 337006
rect 472624 336942 472676 336948
rect 472256 3528 472308 3534
rect 472256 3470 472308 3476
rect 470888 598 471100 626
rect 470888 490 470916 598
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 462 470916 490
rect 471072 480 471100 598
rect 472268 480 472296 3470
rect 472636 3466 472664 336942
rect 560944 336932 560996 336938
rect 560944 336874 560996 336880
rect 497464 336116 497516 336122
rect 497464 336058 497516 336064
rect 480260 335028 480312 335034
rect 480260 334970 480312 334976
rect 476120 332512 476172 332518
rect 476120 332454 476172 332460
rect 474740 329520 474792 329526
rect 474740 329462 474792 329468
rect 474752 3482 474780 329462
rect 476132 16574 476160 332454
rect 477500 327888 477552 327894
rect 477500 327830 477552 327836
rect 477512 16574 477540 327830
rect 480272 16574 480300 334970
rect 483020 334960 483072 334966
rect 483020 334902 483072 334908
rect 481640 332444 481692 332450
rect 481640 332386 481692 332392
rect 476132 16546 476528 16574
rect 477512 16546 478184 16574
rect 480272 16546 480576 16574
rect 472624 3460 472676 3466
rect 472624 3402 472676 3408
rect 473452 3460 473504 3466
rect 473452 3402 473504 3408
rect 474568 3454 474780 3482
rect 475752 3528 475804 3534
rect 475752 3470 475804 3476
rect 473464 480 473492 3402
rect 474568 480 474596 3454
rect 475764 480 475792 3470
rect 476500 490 476528 16546
rect 476776 598 476988 626
rect 476776 490 476804 598
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476500 462 476804 490
rect 476960 480 476988 598
rect 478156 480 478184 16546
rect 479338 3768 479394 3777
rect 479338 3703 479394 3712
rect 479352 480 479380 3703
rect 480548 480 480576 16546
rect 481652 6914 481680 332386
rect 481732 326664 481784 326670
rect 481732 326606 481784 326612
rect 481744 16574 481772 326606
rect 481744 16546 482416 16574
rect 481652 6886 481772 6914
rect 481744 480 481772 6886
rect 482388 490 482416 16546
rect 483032 6914 483060 334902
rect 487160 334892 487212 334898
rect 487160 334834 487212 334840
rect 484400 332376 484452 332382
rect 484400 332318 484452 332324
rect 483664 322312 483716 322318
rect 483664 322254 483716 322260
rect 483676 16574 483704 322254
rect 484412 16574 484440 332318
rect 485780 326596 485832 326602
rect 485780 326538 485832 326544
rect 485792 16574 485820 326538
rect 483676 16546 483796 16574
rect 484412 16546 484808 16574
rect 485792 16546 486464 16574
rect 483032 6886 483704 6914
rect 483676 3346 483704 6886
rect 483768 3466 483796 16546
rect 483756 3460 483808 3466
rect 483756 3402 483808 3408
rect 483676 3318 484072 3346
rect 482664 598 482876 626
rect 482664 490 482692 598
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 462 482692 490
rect 482848 480 482876 598
rect 484044 480 484072 3318
rect 484780 490 484808 16546
rect 485056 598 485268 626
rect 485056 490 485084 598
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 484780 462 485084 490
rect 485240 480 485268 598
rect 486436 480 486464 16546
rect 487172 490 487200 334834
rect 489920 333736 489972 333742
rect 489920 333678 489972 333684
rect 488540 331084 488592 331090
rect 488540 331026 488592 331032
rect 488552 16574 488580 331026
rect 489932 16574 489960 333678
rect 490564 331016 490616 331022
rect 490564 330958 490616 330964
rect 488552 16546 488856 16574
rect 489932 16546 490512 16574
rect 487448 598 487660 626
rect 487448 490 487476 598
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487172 462 487476 490
rect 487632 480 487660 598
rect 488828 480 488856 16546
rect 489920 9104 489972 9110
rect 489920 9046 489972 9052
rect 489932 480 489960 9046
rect 490484 626 490512 16546
rect 490576 3262 490604 330958
rect 492680 326528 492732 326534
rect 492680 326470 492732 326476
rect 492692 16574 492720 326470
rect 496820 325168 496872 325174
rect 496820 325110 496872 325116
rect 496832 16574 496860 325110
rect 492692 16546 493088 16574
rect 496832 16546 497136 16574
rect 490564 3256 490616 3262
rect 490564 3198 490616 3204
rect 492312 3256 492364 3262
rect 492312 3198 492364 3204
rect 490484 598 490696 626
rect 490668 490 490696 598
rect 490944 598 491156 626
rect 490944 490 490972 598
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490668 462 490972 490
rect 491128 480 491156 598
rect 492324 480 492352 3198
rect 493060 490 493088 16546
rect 495900 5092 495952 5098
rect 495900 5034 495952 5040
rect 494704 5024 494756 5030
rect 494704 4966 494756 4972
rect 493336 598 493548 626
rect 493336 490 493364 598
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493060 462 493364 490
rect 493520 480 493548 598
rect 494716 480 494744 4966
rect 495912 480 495940 5034
rect 497108 480 497136 16546
rect 497476 4214 497504 336058
rect 522304 336048 522356 336054
rect 522304 335990 522356 335996
rect 500960 334824 501012 334830
rect 500960 334766 501012 334772
rect 499672 332308 499724 332314
rect 499672 332250 499724 332256
rect 499580 323672 499632 323678
rect 499580 323614 499632 323620
rect 499592 4214 499620 323614
rect 497464 4208 497516 4214
rect 497464 4150 497516 4156
rect 498200 4208 498252 4214
rect 498200 4150 498252 4156
rect 499580 4208 499632 4214
rect 499580 4150 499632 4156
rect 498212 480 498240 4150
rect 499684 4026 499712 332250
rect 500972 16574 501000 334766
rect 514760 334756 514812 334762
rect 514760 334698 514812 334704
rect 507860 333668 507912 333674
rect 507860 333610 507912 333616
rect 506480 333600 506532 333606
rect 506480 333542 506532 333548
rect 502340 330948 502392 330954
rect 502340 330890 502392 330896
rect 502352 16574 502380 330890
rect 503720 327820 503772 327826
rect 503720 327762 503772 327768
rect 500972 16546 501368 16574
rect 502352 16546 503024 16574
rect 500592 4208 500644 4214
rect 500592 4150 500644 4156
rect 499408 3998 499712 4026
rect 499408 480 499436 3998
rect 500604 480 500632 4150
rect 501340 490 501368 16546
rect 501616 598 501828 626
rect 501616 490 501644 598
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501340 462 501644 490
rect 501800 480 501828 598
rect 502996 480 503024 16546
rect 503732 490 503760 327762
rect 505376 4956 505428 4962
rect 505376 4898 505428 4904
rect 504008 598 504220 626
rect 504008 490 504036 598
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 462 504036 490
rect 504192 480 504220 598
rect 505388 480 505416 4898
rect 506492 480 506520 333542
rect 506572 326460 506624 326466
rect 506572 326402 506624 326408
rect 506584 16574 506612 326402
rect 507872 16574 507900 333610
rect 510712 332240 510764 332246
rect 510712 332182 510764 332188
rect 510620 325100 510672 325106
rect 510620 325042 510672 325048
rect 506584 16546 507256 16574
rect 507872 16546 508912 16574
rect 507228 490 507256 16546
rect 507504 598 507716 626
rect 507504 490 507532 598
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 462 507532 490
rect 507688 480 507716 598
rect 508884 480 508912 16546
rect 510068 3528 510120 3534
rect 510068 3470 510120 3476
rect 510080 480 510108 3470
rect 510632 3346 510660 325042
rect 510724 3534 510752 332182
rect 512644 330880 512696 330886
rect 512644 330822 512696 330828
rect 512000 289128 512052 289134
rect 512000 289070 512052 289076
rect 510712 3528 510764 3534
rect 510712 3470 510764 3476
rect 510632 3318 511304 3346
rect 511276 480 511304 3318
rect 512012 490 512040 289070
rect 512656 3534 512684 330822
rect 514772 3602 514800 334698
rect 520280 332104 520332 332110
rect 520280 332046 520332 332052
rect 517520 329452 517572 329458
rect 517520 329394 517572 329400
rect 514852 323604 514904 323610
rect 514852 323546 514904 323552
rect 514760 3596 514812 3602
rect 514760 3538 514812 3544
rect 512644 3528 512696 3534
rect 512644 3470 512696 3476
rect 513564 3528 513616 3534
rect 514864 3482 514892 323546
rect 515956 3596 516008 3602
rect 515956 3538 516008 3544
rect 513564 3470 513616 3476
rect 512288 598 512500 626
rect 512288 490 512316 598
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512012 462 512316 490
rect 512472 480 512500 598
rect 513576 480 513604 3470
rect 514772 3454 514892 3482
rect 514772 480 514800 3454
rect 515968 480 515996 3538
rect 517532 3482 517560 329394
rect 519544 326392 519596 326398
rect 519544 326334 519596 326340
rect 518900 177336 518952 177342
rect 518900 177278 518952 177284
rect 518912 16574 518940 177278
rect 518912 16546 519492 16574
rect 517888 13184 517940 13190
rect 517888 13126 517940 13132
rect 517164 3454 517560 3482
rect 517164 480 517192 3454
rect 517900 490 517928 13126
rect 519464 3346 519492 16546
rect 519556 3534 519584 326334
rect 519544 3528 519596 3534
rect 519544 3470 519596 3476
rect 519464 3318 519584 3346
rect 518176 598 518388 626
rect 518176 490 518204 598
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 462 518204 490
rect 518360 480 518388 598
rect 519556 480 519584 3318
rect 520292 490 520320 332046
rect 522316 4214 522344 335990
rect 543738 335064 543794 335073
rect 543738 334999 543794 335008
rect 532700 334688 532752 334694
rect 532700 334630 532752 334636
rect 529940 333532 529992 333538
rect 529940 333474 529992 333480
rect 524512 333464 524564 333470
rect 524512 333406 524564 333412
rect 524420 325032 524472 325038
rect 524420 324974 524472 324980
rect 522304 4208 522356 4214
rect 522304 4150 522356 4156
rect 523040 4208 523092 4214
rect 523040 4150 523092 4156
rect 521844 3528 521896 3534
rect 521844 3470 521896 3476
rect 520568 598 520780 626
rect 520568 490 520596 598
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520292 462 520596 490
rect 520752 480 520780 598
rect 521856 480 521884 3470
rect 523052 480 523080 4150
rect 524432 3602 524460 324974
rect 524420 3596 524472 3602
rect 524420 3538 524472 3544
rect 524524 3482 524552 333406
rect 525800 332172 525852 332178
rect 525800 332114 525852 332120
rect 525812 16574 525840 332114
rect 528652 330744 528704 330750
rect 528652 330686 528704 330692
rect 528560 322244 528612 322250
rect 528560 322186 528612 322192
rect 525812 16546 526208 16574
rect 525432 3596 525484 3602
rect 525432 3538 525484 3544
rect 524248 3454 524552 3482
rect 524248 480 524276 3454
rect 525444 480 525472 3538
rect 526180 490 526208 16546
rect 527824 3052 527876 3058
rect 527824 2994 527876 3000
rect 526456 598 526668 626
rect 526456 490 526484 598
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526180 462 526484 490
rect 526640 480 526668 598
rect 527836 480 527864 2994
rect 528572 490 528600 322186
rect 528664 3058 528692 330686
rect 529952 16574 529980 333474
rect 530584 329384 530636 329390
rect 530584 329326 530636 329332
rect 529952 16546 530164 16574
rect 528652 3052 528704 3058
rect 528652 2994 528704 3000
rect 528848 598 529060 626
rect 528848 490 528876 598
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528572 462 528876 490
rect 529032 480 529060 598
rect 530136 480 530164 16546
rect 530596 3534 530624 329326
rect 532712 16574 532740 334630
rect 535460 334620 535512 334626
rect 535460 334562 535512 334568
rect 532712 16546 533752 16574
rect 532516 4888 532568 4894
rect 532516 4830 532568 4836
rect 530584 3528 530636 3534
rect 530584 3470 530636 3476
rect 531320 3528 531372 3534
rect 531320 3470 531372 3476
rect 531332 480 531360 3470
rect 532528 480 532556 4830
rect 533724 480 533752 16546
rect 535472 3534 535500 334562
rect 542452 333396 542504 333402
rect 542452 333338 542504 333344
rect 539692 332036 539744 332042
rect 539692 331978 539744 331984
rect 538220 331968 538272 331974
rect 538220 331910 538272 331916
rect 536840 330812 536892 330818
rect 536840 330754 536892 330760
rect 536852 16574 536880 330754
rect 538232 16574 538260 331910
rect 539704 16574 539732 331978
rect 542360 324964 542412 324970
rect 542360 324906 542412 324912
rect 536852 16546 537248 16574
rect 538232 16546 538444 16574
rect 539704 16546 540376 16574
rect 534908 3528 534960 3534
rect 534908 3470 534960 3476
rect 535460 3528 535512 3534
rect 535460 3470 535512 3476
rect 534920 480 534948 3470
rect 536104 3392 536156 3398
rect 536104 3334 536156 3340
rect 536116 480 536144 3334
rect 537220 480 537248 16546
rect 538416 480 538444 16546
rect 539600 3664 539652 3670
rect 539600 3606 539652 3612
rect 539612 480 539640 3606
rect 540348 490 540376 16546
rect 541992 3528 542044 3534
rect 541992 3470 542044 3476
rect 540624 598 540836 626
rect 540624 490 540652 598
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540348 462 540652 490
rect 540808 480 540836 598
rect 542004 480 542032 3470
rect 542372 626 542400 324906
rect 542464 3534 542492 333338
rect 543752 16574 543780 334999
rect 554778 334928 554834 334937
rect 554778 334863 554834 334872
rect 547880 333328 547932 333334
rect 547880 333270 547932 333276
rect 546500 330676 546552 330682
rect 546500 330618 546552 330624
rect 543752 16546 544424 16574
rect 542452 3528 542504 3534
rect 542452 3470 542504 3476
rect 542372 598 542768 626
rect 542740 490 542768 598
rect 543016 598 543228 626
rect 543016 490 543044 598
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542740 462 543044 490
rect 543200 480 543228 598
rect 544396 480 544424 16546
rect 546512 3534 546540 330618
rect 546684 3800 546736 3806
rect 546684 3742 546736 3748
rect 545488 3528 545540 3534
rect 545488 3470 545540 3476
rect 546500 3528 546552 3534
rect 546500 3470 546552 3476
rect 545500 480 545528 3470
rect 546696 480 546724 3742
rect 547892 480 547920 333270
rect 547972 331900 548024 331906
rect 547972 331842 548024 331848
rect 547984 16574 548012 331842
rect 551284 329248 551336 329254
rect 551284 329190 551336 329196
rect 550640 17264 550692 17270
rect 550640 17206 550692 17212
rect 550652 16574 550680 17206
rect 547984 16546 548656 16574
rect 550652 16546 551048 16574
rect 548628 490 548656 16546
rect 550272 3868 550324 3874
rect 550272 3810 550324 3816
rect 548904 598 549116 626
rect 548904 490 548932 598
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 548628 462 548932 490
rect 549088 480 549116 598
rect 550284 480 550312 3810
rect 551020 490 551048 16546
rect 551296 3534 551324 329190
rect 554792 16574 554820 334863
rect 557538 334792 557594 334801
rect 557538 334727 557594 334736
rect 556160 329180 556212 329186
rect 556160 329122 556212 329128
rect 554792 16546 555004 16574
rect 551284 3528 551336 3534
rect 551284 3470 551336 3476
rect 552664 3528 552716 3534
rect 552664 3470 552716 3476
rect 551296 598 551508 626
rect 551296 490 551324 598
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551020 462 551324 490
rect 551480 480 551508 598
rect 552676 480 552704 3470
rect 553768 3460 553820 3466
rect 553768 3402 553820 3408
rect 553780 480 553808 3402
rect 554976 480 555004 16546
rect 556172 480 556200 329122
rect 557552 16574 557580 334727
rect 560300 327752 560352 327758
rect 560300 327694 560352 327700
rect 557552 16546 558592 16574
rect 556896 13116 556948 13122
rect 556896 13058 556948 13064
rect 556908 490 556936 13058
rect 557184 598 557396 626
rect 557184 490 557212 598
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 556908 462 557212 490
rect 557368 480 557396 598
rect 558564 480 558592 16546
rect 560312 3534 560340 327694
rect 560852 4140 560904 4146
rect 560852 4082 560904 4088
rect 559748 3528 559800 3534
rect 559748 3470 559800 3476
rect 560300 3528 560352 3534
rect 560300 3470 560352 3476
rect 559760 480 559788 3470
rect 560864 480 560892 4082
rect 560956 3194 560984 336874
rect 574100 336864 574152 336870
rect 574100 336806 574152 336812
rect 566462 334656 566518 334665
rect 566462 334591 566518 334600
rect 564532 330608 564584 330614
rect 564532 330550 564584 330556
rect 561680 329316 561732 329322
rect 561680 329258 561732 329264
rect 561692 16574 561720 329258
rect 564544 16574 564572 330550
rect 565820 330540 565872 330546
rect 565820 330482 565872 330488
rect 561692 16546 562088 16574
rect 564544 16546 565216 16574
rect 560944 3188 560996 3194
rect 560944 3130 560996 3136
rect 562060 480 562088 16546
rect 564440 3936 564492 3942
rect 564440 3878 564492 3884
rect 563244 3188 563296 3194
rect 563244 3130 563296 3136
rect 563256 480 563284 3130
rect 564452 480 564480 3878
rect 565188 490 565216 16546
rect 565832 6914 565860 330482
rect 566476 16574 566504 334591
rect 568580 333260 568632 333266
rect 568580 333202 568632 333208
rect 568592 16574 568620 333202
rect 569960 329112 570012 329118
rect 569960 329054 570012 329060
rect 569972 16574 570000 329054
rect 574112 16574 574140 336806
rect 580172 325644 580224 325650
rect 580172 325586 580224 325592
rect 580184 325281 580212 325586
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 583116 165912 583168 165918
rect 583114 165880 583116 165889
rect 583168 165880 583170 165889
rect 583114 165815 583170 165824
rect 583024 152720 583076 152726
rect 583022 152688 583024 152697
rect 583076 152688 583078 152697
rect 583022 152623 583078 152632
rect 582840 126064 582892 126070
rect 582838 126032 582840 126041
rect 582892 126032 582894 126041
rect 582838 125967 582894 125976
rect 582748 112872 582800 112878
rect 582746 112840 582748 112849
rect 582800 112840 582802 112849
rect 582746 112775 582802 112784
rect 582656 99544 582708 99550
rect 582654 99512 582656 99521
rect 582708 99512 582710 99521
rect 582654 99447 582710 99456
rect 582564 86216 582616 86222
rect 582562 86184 582564 86193
rect 582616 86184 582618 86193
rect 582562 86119 582618 86128
rect 582472 73024 582524 73030
rect 582470 72992 582472 73001
rect 582524 72992 582526 73001
rect 582470 72927 582526 72936
rect 582380 46368 582432 46374
rect 582378 46336 582380 46345
rect 582432 46336 582434 46345
rect 582378 46271 582434 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 566476 16546 566596 16574
rect 568592 16546 568712 16574
rect 569972 16546 570368 16574
rect 574112 16546 575152 16574
rect 565832 6886 566504 6914
rect 566476 3346 566504 6886
rect 566568 3466 566596 16546
rect 568028 4004 568080 4010
rect 568028 3946 568080 3952
rect 566556 3460 566608 3466
rect 566556 3402 566608 3408
rect 566476 3318 566872 3346
rect 565464 598 565676 626
rect 565464 490 565492 598
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565188 462 565492 490
rect 565648 480 565676 598
rect 566844 480 566872 3318
rect 568040 480 568068 3946
rect 568684 490 568712 16546
rect 568960 598 569172 626
rect 568960 490 568988 598
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 568684 462 568988 490
rect 569144 480 569172 598
rect 570340 480 570368 16546
rect 573916 9036 573968 9042
rect 573916 8978 573968 8984
rect 571524 4072 571576 4078
rect 571524 4014 571576 4020
rect 571536 480 571564 4014
rect 572720 3460 572772 3466
rect 572720 3402 572772 3408
rect 572732 480 572760 3402
rect 573928 480 573956 8978
rect 575124 480 575152 16546
rect 577412 8968 577464 8974
rect 577412 8910 577464 8916
rect 576308 4820 576360 4826
rect 576308 4762 576360 4768
rect 576320 480 576348 4762
rect 577424 480 577452 8910
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 580998 3632 581054 3641
rect 580998 3567 581054 3576
rect 578608 3256 578660 3262
rect 578608 3198 578660 3204
rect 578620 480 578648 3198
rect 581012 480 581040 3567
rect 582194 3496 582250 3505
rect 582194 3431 582250 3440
rect 582208 480 582236 3431
rect 583390 3360 583446 3369
rect 583390 3295 583446 3304
rect 583404 480 583432 3295
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3146 658144 3202 658200
rect 3330 606056 3386 606112
rect 3146 553832 3202 553888
rect 3238 501744 3294 501800
rect 3330 475632 3386 475688
rect 3238 462576 3294 462632
rect 3146 449520 3202 449576
rect 3146 423544 3202 423600
rect 3054 410488 3110 410544
rect 2962 397468 2964 397488
rect 2964 397468 3016 397488
rect 3016 397468 3018 397488
rect 2962 397432 3018 397468
rect 3514 671200 3570 671256
rect 3606 632032 3662 632088
rect 3698 619112 3754 619168
rect 3790 579944 3846 580000
rect 3882 566888 3938 566944
rect 3974 527856 4030 527912
rect 4066 514800 4122 514856
rect 24766 380296 24822 380352
rect 3422 380160 3478 380216
rect 3146 345344 3202 345400
rect 3054 293120 3110 293176
rect 3330 214920 3386 214976
rect 2778 162832 2834 162888
rect 3606 371320 3662 371376
rect 3514 358400 3570 358456
rect 3514 319232 3570 319288
rect 3514 306176 3570 306232
rect 3514 267144 3570 267200
rect 3514 255176 3570 255232
rect 3514 254088 3570 254144
rect 3514 241032 3570 241088
rect 3514 202816 3570 202872
rect 3514 201864 3570 201920
rect 3514 188808 3570 188864
rect 3514 137944 3570 138000
rect 3514 136720 3570 136776
rect 3422 110608 3478 110664
rect 3146 84632 3202 84688
rect 3422 71576 3478 71632
rect 3330 59200 3386 59256
rect 3330 58520 3386 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3146 32408 3202 32464
rect 3422 19352 3478 19408
rect 3330 6432 3386 6488
rect 6458 3304 6514 3360
rect 25502 336096 25558 336152
rect 14462 335960 14518 336016
rect 15934 3576 15990 3632
rect 14738 3440 14794 3496
rect 20626 3712 20682 3768
rect 177302 336640 177358 336696
rect 173162 336504 173218 336560
rect 130382 336232 130438 336288
rect 180062 336368 180118 336424
rect 272246 380296 272302 380352
rect 272706 380160 272762 380216
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 458088 580226 458144
rect 580170 431568 580226 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 234526 335824 234582 335880
rect 235446 377304 235502 377360
rect 236550 377304 236606 377360
rect 238114 377304 238170 377360
rect 241242 377304 241298 377360
rect 242714 377304 242770 377360
rect 244002 377304 244058 377360
rect 286414 377304 286470 377360
rect 287978 377304 288034 377360
rect 289082 377304 289138 377360
rect 290186 377304 290242 377360
rect 291198 377304 291254 377360
rect 292762 377304 292818 377360
rect 294326 377304 294382 377360
rect 234710 377168 234766 377224
rect 294970 377168 295026 377224
rect 235446 336504 235502 336560
rect 235906 336640 235962 336696
rect 236090 335960 236146 336016
rect 234802 3304 234858 3360
rect 236182 3576 236238 3632
rect 236918 336096 236974 336152
rect 237838 336232 237894 336288
rect 236550 3712 236606 3768
rect 236366 3440 236422 3496
rect 245014 335416 245070 335472
rect 245474 336368 245530 336424
rect 247130 335416 247186 335472
rect 247866 335824 247922 335880
rect 272890 335996 272892 336016
rect 272892 335996 272944 336016
rect 272944 335996 272946 336016
rect 272890 335960 272946 335996
rect 272890 335552 272946 335608
rect 274914 336096 274970 336152
rect 275282 337592 275338 337648
rect 275742 337864 275798 337920
rect 275650 335688 275706 335744
rect 278318 335960 278374 336016
rect 278318 335572 278374 335608
rect 278318 335552 278320 335572
rect 278320 335552 278372 335572
rect 278372 335552 278374 335572
rect 279330 335552 279386 335608
rect 282458 335416 282514 335472
rect 282826 336096 282882 336152
rect 282918 335960 282974 336016
rect 282826 335688 282882 335744
rect 282826 335416 282882 335472
rect 283102 335416 283158 335472
rect 284114 3712 284170 3768
rect 284850 335552 284906 335608
rect 286506 335416 286562 335472
rect 287334 335960 287390 336016
rect 288346 335960 288402 336016
rect 290278 336232 290334 336288
rect 291014 335416 291070 335472
rect 291428 337864 291484 337920
rect 291382 336504 291438 336560
rect 291658 336096 291714 336152
rect 292026 334872 292082 334928
rect 292394 334736 292450 334792
rect 293130 335552 293186 335608
rect 293590 335688 293646 335744
rect 293958 334600 294014 334656
rect 295522 337864 295578 337920
rect 295246 3576 295302 3632
rect 295154 3440 295210 3496
rect 295062 3304 295118 3360
rect 295798 335552 295854 335608
rect 296442 336504 296498 336560
rect 298006 335688 298062 335744
rect 299938 336232 299994 336288
rect 580170 378428 580172 378448
rect 580172 378428 580224 378448
rect 580224 378428 580226 378448
rect 580170 378392 580226 378428
rect 580170 365064 580226 365120
rect 580170 351872 580226 351928
rect 327722 336096 327778 336152
rect 324962 335960 325018 336016
rect 479338 3712 479394 3768
rect 543738 335008 543794 335064
rect 554778 334872 554834 334928
rect 557538 334736 557594 334792
rect 566462 334600 566518 334656
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 580170 258848 580226 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 579986 232328 580042 232384
rect 579802 205672 579858 205728
rect 580170 192480 580226 192536
rect 583114 165860 583116 165880
rect 583116 165860 583168 165880
rect 583168 165860 583170 165880
rect 583114 165824 583170 165860
rect 583022 152668 583024 152688
rect 583024 152668 583076 152688
rect 583076 152668 583078 152688
rect 583022 152632 583078 152668
rect 582838 126012 582840 126032
rect 582840 126012 582892 126032
rect 582892 126012 582894 126032
rect 582838 125976 582894 126012
rect 582746 112820 582748 112840
rect 582748 112820 582800 112840
rect 582800 112820 582802 112840
rect 582746 112784 582802 112820
rect 582654 99492 582656 99512
rect 582656 99492 582708 99512
rect 582708 99492 582710 99512
rect 582654 99456 582710 99492
rect 582562 86164 582564 86184
rect 582564 86164 582616 86184
rect 582616 86164 582618 86184
rect 582562 86128 582618 86164
rect 582470 72972 582472 72992
rect 582472 72972 582524 72992
rect 582524 72972 582526 72992
rect 582470 72936 582526 72972
rect 582378 46316 582380 46336
rect 582380 46316 582432 46336
rect 582432 46316 582434 46336
rect 582378 46280 582434 46316
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 580170 6568 580226 6624
rect 580998 3576 581054 3632
rect 582194 3440 582250 3496
rect 583390 3304 583446 3360
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3141 658202 3207 658205
rect -960 658200 3207 658202
rect -960 658144 3146 658200
rect 3202 658144 3207 658200
rect -960 658142 3207 658144
rect -960 658052 480 658142
rect 3141 658139 3207 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3601 632090 3667 632093
rect -960 632088 3667 632090
rect -960 632032 3606 632088
rect 3662 632032 3667 632088
rect -960 632030 3667 632032
rect -960 631940 480 632030
rect 3601 632027 3667 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3693 619170 3759 619173
rect -960 619168 3759 619170
rect -960 619112 3698 619168
rect 3754 619112 3759 619168
rect -960 619110 3759 619112
rect -960 619020 480 619110
rect 3693 619107 3759 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3325 606114 3391 606117
rect -960 606112 3391 606114
rect -960 606056 3330 606112
rect 3386 606056 3391 606112
rect -960 606054 3391 606056
rect -960 605964 480 606054
rect 3325 606051 3391 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3785 580002 3851 580005
rect -960 580000 3851 580002
rect -960 579944 3790 580000
rect 3846 579944 3851 580000
rect -960 579942 3851 579944
rect -960 579852 480 579942
rect 3785 579939 3851 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3877 566946 3943 566949
rect -960 566944 3943 566946
rect -960 566888 3882 566944
rect 3938 566888 3943 566944
rect -960 566886 3943 566888
rect -960 566796 480 566886
rect 3877 566883 3943 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3141 553890 3207 553893
rect -960 553888 3207 553890
rect -960 553832 3146 553888
rect 3202 553832 3207 553888
rect -960 553830 3207 553832
rect -960 553740 480 553830
rect 3141 553827 3207 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3969 527914 4035 527917
rect -960 527912 4035 527914
rect -960 527856 3974 527912
rect 4030 527856 4035 527912
rect -960 527854 4035 527856
rect -960 527764 480 527854
rect 3969 527851 4035 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 4061 514858 4127 514861
rect -960 514856 4127 514858
rect -960 514800 4066 514856
rect 4122 514800 4127 514856
rect -960 514798 4127 514800
rect -960 514708 480 514798
rect 4061 514795 4127 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3233 501802 3299 501805
rect -960 501800 3299 501802
rect -960 501744 3238 501800
rect 3294 501744 3299 501800
rect -960 501742 3299 501744
rect -960 501652 480 501742
rect 3233 501739 3299 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3325 475690 3391 475693
rect -960 475688 3391 475690
rect -960 475632 3330 475688
rect 3386 475632 3391 475688
rect -960 475630 3391 475632
rect -960 475540 480 475630
rect 3325 475627 3391 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3233 462634 3299 462637
rect -960 462632 3299 462634
rect -960 462576 3238 462632
rect 3294 462576 3299 462632
rect -960 462574 3299 462576
rect -960 462484 480 462574
rect 3233 462571 3299 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3141 423602 3207 423605
rect -960 423600 3207 423602
rect -960 423544 3146 423600
rect 3202 423544 3207 423600
rect -960 423542 3207 423544
rect -960 423452 480 423542
rect 3141 423539 3207 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3049 410546 3115 410549
rect -960 410544 3115 410546
rect -960 410488 3054 410544
rect 3110 410488 3115 410544
rect -960 410486 3115 410488
rect -960 410396 480 410486
rect 3049 410483 3115 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 2957 397490 3023 397493
rect -960 397488 3023 397490
rect -960 397432 2962 397488
rect 3018 397432 3023 397488
rect -960 397430 3023 397432
rect -960 397340 480 397430
rect 2957 397427 3023 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 24761 380354 24827 380357
rect 272241 380354 272307 380357
rect 24761 380352 272307 380354
rect 24761 380296 24766 380352
rect 24822 380296 272246 380352
rect 272302 380296 272307 380352
rect 24761 380294 272307 380296
rect 24761 380291 24827 380294
rect 272241 380291 272307 380294
rect 3417 380218 3483 380221
rect 272701 380218 272767 380221
rect 3417 380216 272767 380218
rect 3417 380160 3422 380216
rect 3478 380160 272706 380216
rect 272762 380160 272767 380216
rect 3417 380158 272767 380160
rect 3417 380155 3483 380158
rect 272701 380155 272767 380158
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 235441 377362 235507 377365
rect 234846 377360 235507 377362
rect 234846 377304 235446 377360
rect 235502 377304 235507 377360
rect 234846 377302 235507 377304
rect 234705 377226 234771 377229
rect 234846 377226 234906 377302
rect 235441 377299 235507 377302
rect 236545 377362 236611 377365
rect 237230 377362 237236 377364
rect 236545 377360 237236 377362
rect 236545 377304 236550 377360
rect 236606 377304 237236 377360
rect 236545 377302 237236 377304
rect 236545 377299 236611 377302
rect 237230 377300 237236 377302
rect 237300 377300 237306 377364
rect 238109 377362 238175 377365
rect 241237 377364 241303 377365
rect 242709 377364 242775 377365
rect 243997 377364 244063 377365
rect 238518 377362 238524 377364
rect 238109 377360 238524 377362
rect 238109 377304 238114 377360
rect 238170 377304 238524 377360
rect 238109 377302 238524 377304
rect 238109 377299 238175 377302
rect 238518 377300 238524 377302
rect 238588 377300 238594 377364
rect 241237 377360 241284 377364
rect 241348 377362 241354 377364
rect 241237 377304 241242 377360
rect 241237 377300 241284 377304
rect 241348 377302 241394 377362
rect 242709 377360 242756 377364
rect 242820 377362 242826 377364
rect 242709 377304 242714 377360
rect 241348 377300 241354 377302
rect 242709 377300 242756 377304
rect 242820 377302 242866 377362
rect 243997 377360 244044 377364
rect 244108 377362 244114 377364
rect 243997 377304 244002 377360
rect 242820 377300 242826 377302
rect 243997 377300 244044 377304
rect 244108 377302 244154 377362
rect 244108 377300 244114 377302
rect 285806 377300 285812 377364
rect 285876 377362 285882 377364
rect 286409 377362 286475 377365
rect 285876 377360 286475 377362
rect 285876 377304 286414 377360
rect 286470 377304 286475 377360
rect 285876 377302 286475 377304
rect 285876 377300 285882 377302
rect 241237 377299 241303 377300
rect 242709 377299 242775 377300
rect 243997 377299 244063 377300
rect 286409 377299 286475 377302
rect 287094 377300 287100 377364
rect 287164 377362 287170 377364
rect 287973 377362 288039 377365
rect 287164 377360 288039 377362
rect 287164 377304 287978 377360
rect 288034 377304 288039 377360
rect 287164 377302 288039 377304
rect 287164 377300 287170 377302
rect 287973 377299 288039 377302
rect 288382 377300 288388 377364
rect 288452 377362 288458 377364
rect 289077 377362 289143 377365
rect 288452 377360 289143 377362
rect 288452 377304 289082 377360
rect 289138 377304 289143 377360
rect 288452 377302 289143 377304
rect 288452 377300 288458 377302
rect 289077 377299 289143 377302
rect 290181 377362 290247 377365
rect 291193 377364 291259 377365
rect 290590 377362 290596 377364
rect 290181 377360 290596 377362
rect 290181 377304 290186 377360
rect 290242 377304 290596 377360
rect 290181 377302 290596 377304
rect 290181 377299 290247 377302
rect 290590 377300 290596 377302
rect 290660 377300 290666 377364
rect 291142 377362 291148 377364
rect 291102 377302 291148 377362
rect 291212 377360 291259 377364
rect 291254 377304 291259 377360
rect 291142 377300 291148 377302
rect 291212 377300 291259 377304
rect 292614 377300 292620 377364
rect 292684 377362 292690 377364
rect 292757 377362 292823 377365
rect 292684 377360 292823 377362
rect 292684 377304 292762 377360
rect 292818 377304 292823 377360
rect 292684 377302 292823 377304
rect 292684 377300 292690 377302
rect 291193 377299 291259 377300
rect 292757 377299 292823 377302
rect 294321 377362 294387 377365
rect 294321 377360 294522 377362
rect 294321 377304 294326 377360
rect 294382 377304 294522 377360
rect 294321 377302 294522 377304
rect 294321 377299 294387 377302
rect 234705 377224 234906 377226
rect 234705 377168 234710 377224
rect 234766 377168 234906 377224
rect 234705 377166 234906 377168
rect 294462 377226 294522 377302
rect 294965 377226 295031 377229
rect 294462 377224 295031 377226
rect 294462 377168 294970 377224
rect 295026 377168 295031 377224
rect 294462 377166 295031 377168
rect 234705 377163 234771 377166
rect 294965 377163 295031 377166
rect -960 371378 480 371468
rect 3601 371378 3667 371381
rect -960 371376 3667 371378
rect -960 371320 3606 371376
rect 3662 371320 3667 371376
rect -960 371318 3667 371320
rect -960 371228 480 371318
rect 3601 371315 3667 371318
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3509 358458 3575 358461
rect -960 358456 3575 358458
rect -960 358400 3514 358456
rect 3570 358400 3575 358456
rect -960 358398 3575 358400
rect -960 358308 480 358398
rect 3509 358395 3575 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3141 345402 3207 345405
rect -960 345400 3207 345402
rect -960 345344 3146 345400
rect 3202 345344 3207 345400
rect -960 345342 3207 345344
rect -960 345252 480 345342
rect 3141 345339 3207 345342
rect 583520 338452 584960 338692
rect 275737 337922 275803 337925
rect 275510 337920 275803 337922
rect 275510 337864 275742 337920
rect 275798 337864 275803 337920
rect 275510 337862 275803 337864
rect 275277 337650 275343 337653
rect 275510 337650 275570 337862
rect 275737 337859 275803 337862
rect 291423 337922 291489 337925
rect 295517 337922 295583 337925
rect 291423 337920 295583 337922
rect 291423 337864 291428 337920
rect 291484 337864 295522 337920
rect 295578 337864 295583 337920
rect 291423 337862 295583 337864
rect 291423 337859 291489 337862
rect 295517 337859 295583 337862
rect 275277 337648 275570 337650
rect 275277 337592 275282 337648
rect 275338 337592 275570 337648
rect 275277 337590 275570 337592
rect 275277 337587 275343 337590
rect 177297 336698 177363 336701
rect 235901 336698 235967 336701
rect 177297 336696 235967 336698
rect 177297 336640 177302 336696
rect 177358 336640 235906 336696
rect 235962 336640 235967 336696
rect 177297 336638 235967 336640
rect 177297 336635 177363 336638
rect 235901 336635 235967 336638
rect 173157 336562 173223 336565
rect 235441 336562 235507 336565
rect 173157 336560 235507 336562
rect 173157 336504 173162 336560
rect 173218 336504 235446 336560
rect 235502 336504 235507 336560
rect 173157 336502 235507 336504
rect 173157 336499 173223 336502
rect 235441 336499 235507 336502
rect 291377 336562 291443 336565
rect 296437 336562 296503 336565
rect 291377 336560 296503 336562
rect 291377 336504 291382 336560
rect 291438 336504 296442 336560
rect 296498 336504 296503 336560
rect 291377 336502 296503 336504
rect 291377 336499 291443 336502
rect 296437 336499 296503 336502
rect 180057 336426 180123 336429
rect 245469 336426 245535 336429
rect 180057 336424 245535 336426
rect 180057 336368 180062 336424
rect 180118 336368 245474 336424
rect 245530 336368 245535 336424
rect 180057 336366 245535 336368
rect 180057 336363 180123 336366
rect 245469 336363 245535 336366
rect 130377 336290 130443 336293
rect 237833 336290 237899 336293
rect 130377 336288 237899 336290
rect 130377 336232 130382 336288
rect 130438 336232 237838 336288
rect 237894 336232 237899 336288
rect 130377 336230 237899 336232
rect 130377 336227 130443 336230
rect 237833 336227 237899 336230
rect 290273 336290 290339 336293
rect 299933 336290 299999 336293
rect 290273 336288 299999 336290
rect 290273 336232 290278 336288
rect 290334 336232 299938 336288
rect 299994 336232 299999 336288
rect 290273 336230 299999 336232
rect 290273 336227 290339 336230
rect 299933 336227 299999 336230
rect 25497 336154 25563 336157
rect 236913 336154 236979 336157
rect 25497 336152 236979 336154
rect 25497 336096 25502 336152
rect 25558 336096 236918 336152
rect 236974 336096 236979 336152
rect 25497 336094 236979 336096
rect 25497 336091 25563 336094
rect 236913 336091 236979 336094
rect 274909 336154 274975 336157
rect 282821 336154 282887 336157
rect 274909 336152 282887 336154
rect 274909 336096 274914 336152
rect 274970 336096 282826 336152
rect 282882 336096 282887 336152
rect 274909 336094 282887 336096
rect 274909 336091 274975 336094
rect 282821 336091 282887 336094
rect 291653 336154 291719 336157
rect 327717 336154 327783 336157
rect 291653 336152 327783 336154
rect 291653 336096 291658 336152
rect 291714 336096 327722 336152
rect 327778 336096 327783 336152
rect 291653 336094 327783 336096
rect 291653 336091 291719 336094
rect 327717 336091 327783 336094
rect 14457 336018 14523 336021
rect 236085 336018 236151 336021
rect 14457 336016 236151 336018
rect 14457 335960 14462 336016
rect 14518 335960 236090 336016
rect 236146 335960 236151 336016
rect 14457 335958 236151 335960
rect 14457 335955 14523 335958
rect 236085 335955 236151 335958
rect 272885 336018 272951 336021
rect 278313 336018 278379 336021
rect 272885 336016 278379 336018
rect 272885 335960 272890 336016
rect 272946 335960 278318 336016
rect 278374 335960 278379 336016
rect 272885 335958 278379 335960
rect 272885 335955 272951 335958
rect 278313 335955 278379 335958
rect 282913 336018 282979 336021
rect 287329 336018 287395 336021
rect 282913 336016 287395 336018
rect 282913 335960 282918 336016
rect 282974 335960 287334 336016
rect 287390 335960 287395 336016
rect 282913 335958 287395 335960
rect 282913 335955 282979 335958
rect 287329 335955 287395 335958
rect 288341 336018 288407 336021
rect 324957 336018 325023 336021
rect 288341 336016 325023 336018
rect 288341 335960 288346 336016
rect 288402 335960 324962 336016
rect 325018 335960 325023 336016
rect 288341 335958 325023 335960
rect 288341 335955 288407 335958
rect 324957 335955 325023 335958
rect 234521 335882 234587 335885
rect 247861 335882 247927 335885
rect 234521 335880 247927 335882
rect 234521 335824 234526 335880
rect 234582 335824 247866 335880
rect 247922 335824 247927 335880
rect 234521 335822 247927 335824
rect 234521 335819 234587 335822
rect 247861 335819 247927 335822
rect 275645 335746 275711 335749
rect 282821 335746 282887 335749
rect 275645 335744 282887 335746
rect 275645 335688 275650 335744
rect 275706 335688 282826 335744
rect 282882 335688 282887 335744
rect 275645 335686 282887 335688
rect 275645 335683 275711 335686
rect 282821 335683 282887 335686
rect 293585 335746 293651 335749
rect 298001 335746 298067 335749
rect 293585 335744 298067 335746
rect 293585 335688 293590 335744
rect 293646 335688 298006 335744
rect 298062 335688 298067 335744
rect 293585 335686 298067 335688
rect 293585 335683 293651 335686
rect 298001 335683 298067 335686
rect 272885 335610 272951 335613
rect 278313 335610 278379 335613
rect 272885 335608 278379 335610
rect 272885 335552 272890 335608
rect 272946 335552 278318 335608
rect 278374 335552 278379 335608
rect 272885 335550 278379 335552
rect 272885 335547 272951 335550
rect 278313 335547 278379 335550
rect 279325 335610 279391 335613
rect 284845 335610 284911 335613
rect 279325 335608 284911 335610
rect 279325 335552 279330 335608
rect 279386 335552 284850 335608
rect 284906 335552 284911 335608
rect 279325 335550 284911 335552
rect 279325 335547 279391 335550
rect 284845 335547 284911 335550
rect 293125 335610 293191 335613
rect 295793 335610 295859 335613
rect 293125 335608 295859 335610
rect 293125 335552 293130 335608
rect 293186 335552 295798 335608
rect 295854 335552 295859 335608
rect 293125 335550 295859 335552
rect 293125 335547 293191 335550
rect 295793 335547 295859 335550
rect 245009 335474 245075 335477
rect 247125 335474 247191 335477
rect 245009 335472 247191 335474
rect 245009 335416 245014 335472
rect 245070 335416 247130 335472
rect 247186 335416 247191 335472
rect 245009 335414 247191 335416
rect 245009 335411 245075 335414
rect 247125 335411 247191 335414
rect 282453 335474 282519 335477
rect 282821 335474 282887 335477
rect 282453 335472 282887 335474
rect 282453 335416 282458 335472
rect 282514 335416 282826 335472
rect 282882 335416 282887 335472
rect 282453 335414 282887 335416
rect 282453 335411 282519 335414
rect 282821 335411 282887 335414
rect 283097 335474 283163 335477
rect 286501 335474 286567 335477
rect 283097 335472 286567 335474
rect 283097 335416 283102 335472
rect 283158 335416 286506 335472
rect 286562 335416 286567 335472
rect 283097 335414 286567 335416
rect 283097 335411 283163 335414
rect 286501 335411 286567 335414
rect 291009 335474 291075 335477
rect 291009 335472 297466 335474
rect 291009 335416 291014 335472
rect 291070 335416 297466 335472
rect 291009 335414 297466 335416
rect 291009 335411 291075 335414
rect 297406 335338 297466 335414
rect 297406 335278 302250 335338
rect 302190 335066 302250 335278
rect 543733 335066 543799 335069
rect 302190 335064 543799 335066
rect 302190 335008 543738 335064
rect 543794 335008 543799 335064
rect 302190 335006 543799 335008
rect 543733 335003 543799 335006
rect 292021 334930 292087 334933
rect 554773 334930 554839 334933
rect 292021 334928 554839 334930
rect 292021 334872 292026 334928
rect 292082 334872 554778 334928
rect 554834 334872 554839 334928
rect 292021 334870 554839 334872
rect 292021 334867 292087 334870
rect 554773 334867 554839 334870
rect 292389 334794 292455 334797
rect 557533 334794 557599 334797
rect 292389 334792 557599 334794
rect 292389 334736 292394 334792
rect 292450 334736 557538 334792
rect 557594 334736 557599 334792
rect 292389 334734 557599 334736
rect 292389 334731 292455 334734
rect 557533 334731 557599 334734
rect 293953 334658 294019 334661
rect 566457 334658 566523 334661
rect 293953 334656 566523 334658
rect 293953 334600 293958 334656
rect 294014 334600 566462 334656
rect 566518 334600 566523 334656
rect 293953 334598 566523 334600
rect 293953 334595 294019 334598
rect 566457 334595 566523 334598
rect -960 332196 480 332436
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3509 319290 3575 319293
rect -960 319288 3575 319290
rect -960 319232 3514 319288
rect 3570 319232 3575 319288
rect -960 319230 3575 319232
rect -960 319140 480 319230
rect 3509 319227 3575 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3509 306234 3575 306237
rect -960 306232 3575 306234
rect -960 306176 3514 306232
rect 3570 306176 3575 306232
rect -960 306174 3575 306176
rect -960 306084 480 306174
rect 3509 306171 3575 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3049 293178 3115 293181
rect -960 293176 3115 293178
rect -960 293120 3054 293176
rect 3110 293120 3115 293176
rect -960 293118 3115 293120
rect -960 293028 480 293118
rect 3049 293115 3115 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3509 267202 3575 267205
rect -960 267200 3575 267202
rect -960 267144 3514 267200
rect 3570 267144 3575 267200
rect -960 267142 3575 267144
rect -960 267052 480 267142
rect 3509 267139 3575 267142
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect 3509 255234 3575 255237
rect 285806 255234 285812 255236
rect 3509 255232 285812 255234
rect 3509 255176 3514 255232
rect 3570 255176 285812 255232
rect 3509 255174 285812 255176
rect 3509 255171 3575 255174
rect 285806 255172 285812 255174
rect 285876 255172 285882 255236
rect -960 254146 480 254236
rect 3509 254146 3575 254149
rect -960 254144 3575 254146
rect -960 254088 3514 254144
rect 3570 254088 3575 254144
rect -960 254086 3575 254088
rect -960 253996 480 254086
rect 3509 254083 3575 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 583520 219058 584960 219148
rect 583342 218998 584960 219058
rect 583342 218922 583402 218998
rect 583520 218922 584960 218998
rect 583342 218908 584960 218922
rect 583342 218862 583586 218908
rect 244038 218044 244044 218108
rect 244108 218106 244114 218108
rect 583526 218106 583586 218862
rect 244108 218046 583586 218106
rect 244108 218044 244114 218046
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect 3509 202874 3575 202877
rect 287094 202874 287100 202876
rect 3509 202872 287100 202874
rect 3509 202816 3514 202872
rect 3570 202816 287100 202872
rect 3509 202814 287100 202816
rect 3509 202811 3575 202814
rect 287094 202812 287100 202814
rect 287164 202812 287170 202876
rect -960 201922 480 202012
rect 3509 201922 3575 201925
rect -960 201920 3575 201922
rect -960 201864 3514 201920
rect 3570 201864 3575 201920
rect -960 201862 3575 201864
rect -960 201772 480 201862
rect 3509 201859 3575 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 583520 179210 584960 179300
rect 583342 179150 584960 179210
rect 583342 179074 583402 179150
rect 583520 179074 584960 179150
rect 583342 179060 584960 179074
rect 583342 179014 583586 179060
rect 242750 178060 242756 178124
rect 242820 178122 242826 178124
rect 583526 178122 583586 179014
rect 242820 178062 583586 178122
rect 242820 178060 242826 178062
rect -960 175796 480 176036
rect 583109 165882 583175 165885
rect 583520 165882 584960 165972
rect 583109 165880 584960 165882
rect 583109 165824 583114 165880
rect 583170 165824 584960 165880
rect 583109 165822 584960 165824
rect 583109 165819 583175 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 2773 162890 2839 162893
rect -960 162888 2839 162890
rect -960 162832 2778 162888
rect 2834 162832 2839 162888
rect -960 162830 2839 162832
rect -960 162740 480 162830
rect 2773 162827 2839 162830
rect 583017 152690 583083 152693
rect 583520 152690 584960 152780
rect 583017 152688 584960 152690
rect 583017 152632 583022 152688
rect 583078 152632 584960 152688
rect 583017 152630 584960 152632
rect 583017 152627 583083 152630
rect 583520 152540 584960 152630
rect 290590 150378 290596 150380
rect 430 150318 290596 150378
rect 430 150106 490 150318
rect 290590 150316 290596 150318
rect 290660 150316 290666 150380
rect 430 150046 674 150106
rect -960 149834 480 149924
rect 614 149834 674 150046
rect -960 149774 674 149834
rect -960 149684 480 149774
rect 583520 139362 584960 139452
rect 583342 139302 584960 139362
rect 583342 139226 583402 139302
rect 583520 139226 584960 139302
rect 583342 139212 584960 139226
rect 583342 139166 583586 139212
rect 241278 138076 241284 138140
rect 241348 138138 241354 138140
rect 583526 138138 583586 139166
rect 241348 138078 583586 138138
rect 241348 138076 241354 138078
rect 3509 138002 3575 138005
rect 288382 138002 288388 138004
rect 3509 138000 288388 138002
rect 3509 137944 3514 138000
rect 3570 137944 288388 138000
rect 3509 137942 288388 137944
rect 3509 137939 3575 137942
rect 288382 137940 288388 137942
rect 288452 137940 288458 138004
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 582833 126034 582899 126037
rect 583520 126034 584960 126124
rect 582833 126032 584960 126034
rect 582833 125976 582838 126032
rect 582894 125976 584960 126032
rect 582833 125974 584960 125976
rect 582833 125971 582899 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 582741 112842 582807 112845
rect 583520 112842 584960 112932
rect 582741 112840 584960 112842
rect 582741 112784 582746 112840
rect 582802 112784 584960 112840
rect 582741 112782 584960 112784
rect 582741 112779 582807 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 582649 99514 582715 99517
rect 583520 99514 584960 99604
rect 582649 99512 584960 99514
rect 582649 99456 582654 99512
rect 582710 99456 584960 99512
rect 582649 99454 584960 99456
rect 582649 99451 582715 99454
rect 583520 99364 584960 99454
rect 291142 97882 291148 97884
rect 6870 97822 291148 97882
rect -960 97610 480 97700
rect 6870 97610 6930 97822
rect 291142 97820 291148 97822
rect 291212 97820 291218 97884
rect -960 97550 6930 97610
rect -960 97460 480 97550
rect 582557 86186 582623 86189
rect 583520 86186 584960 86276
rect 582557 86184 584960 86186
rect 582557 86128 582562 86184
rect 582618 86128 584960 86184
rect 582557 86126 584960 86128
rect 582557 86123 582623 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 582465 72994 582531 72997
rect 583520 72994 584960 73084
rect 582465 72992 584960 72994
rect 582465 72936 582470 72992
rect 582526 72936 584960 72992
rect 582465 72934 584960 72936
rect 582465 72931 582531 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 583520 59666 584960 59756
rect 567150 59606 584960 59666
rect 238518 59332 238524 59396
rect 238588 59394 238594 59396
rect 567150 59394 567210 59606
rect 583520 59516 584960 59606
rect 238588 59334 567210 59394
rect 238588 59332 238594 59334
rect 3325 59258 3391 59261
rect 292614 59258 292620 59260
rect 3325 59256 292620 59258
rect 3325 59200 3330 59256
rect 3386 59200 292620 59256
rect 3325 59198 292620 59200
rect 3325 59195 3391 59198
rect 292614 59196 292620 59198
rect 292684 59196 292690 59260
rect -960 58578 480 58668
rect 3325 58578 3391 58581
rect -960 58576 3391 58578
rect -960 58520 3330 58576
rect 3386 58520 3391 58576
rect -960 58518 3391 58520
rect -960 58428 480 58518
rect 3325 58515 3391 58518
rect 582373 46338 582439 46341
rect 583520 46338 584960 46428
rect 582373 46336 584960 46338
rect 582373 46280 582378 46336
rect 582434 46280 584960 46336
rect 582373 46278 584960 46280
rect 582373 46275 582439 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3141 32466 3207 32469
rect -960 32464 3207 32466
rect -960 32408 3146 32464
rect 3202 32408 3207 32464
rect -960 32406 3207 32408
rect -960 32316 480 32406
rect 3141 32403 3207 32406
rect 583520 19818 584960 19908
rect 583342 19758 584960 19818
rect 583342 19682 583402 19758
rect 583520 19682 584960 19758
rect 583342 19668 584960 19682
rect 583342 19622 583586 19668
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 237230 19348 237236 19412
rect 237300 19410 237306 19412
rect 583526 19410 583586 19622
rect 237300 19350 583586 19410
rect 237300 19348 237306 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3325 6490 3391 6493
rect -960 6488 3391 6490
rect -960 6432 3330 6488
rect 3386 6432 3391 6488
rect 583520 6476 584960 6566
rect -960 6430 3391 6432
rect -960 6340 480 6430
rect 3325 6427 3391 6430
rect 20621 3770 20687 3773
rect 236545 3770 236611 3773
rect 20621 3768 236611 3770
rect 20621 3712 20626 3768
rect 20682 3712 236550 3768
rect 236606 3712 236611 3768
rect 20621 3710 236611 3712
rect 20621 3707 20687 3710
rect 236545 3707 236611 3710
rect 284109 3770 284175 3773
rect 479333 3770 479399 3773
rect 284109 3768 479399 3770
rect 284109 3712 284114 3768
rect 284170 3712 479338 3768
rect 479394 3712 479399 3768
rect 284109 3710 479399 3712
rect 284109 3707 284175 3710
rect 479333 3707 479399 3710
rect 15929 3634 15995 3637
rect 236177 3634 236243 3637
rect 15929 3632 236243 3634
rect 15929 3576 15934 3632
rect 15990 3576 236182 3632
rect 236238 3576 236243 3632
rect 15929 3574 236243 3576
rect 15929 3571 15995 3574
rect 236177 3571 236243 3574
rect 295241 3634 295307 3637
rect 580993 3634 581059 3637
rect 295241 3632 581059 3634
rect 295241 3576 295246 3632
rect 295302 3576 580998 3632
rect 581054 3576 581059 3632
rect 295241 3574 581059 3576
rect 295241 3571 295307 3574
rect 580993 3571 581059 3574
rect 14733 3498 14799 3501
rect 236361 3498 236427 3501
rect 14733 3496 236427 3498
rect 14733 3440 14738 3496
rect 14794 3440 236366 3496
rect 236422 3440 236427 3496
rect 14733 3438 236427 3440
rect 14733 3435 14799 3438
rect 236361 3435 236427 3438
rect 295149 3498 295215 3501
rect 582189 3498 582255 3501
rect 295149 3496 582255 3498
rect 295149 3440 295154 3496
rect 295210 3440 582194 3496
rect 582250 3440 582255 3496
rect 295149 3438 582255 3440
rect 295149 3435 295215 3438
rect 582189 3435 582255 3438
rect 6453 3362 6519 3365
rect 234797 3362 234863 3365
rect 6453 3360 234863 3362
rect 6453 3304 6458 3360
rect 6514 3304 234802 3360
rect 234858 3304 234863 3360
rect 6453 3302 234863 3304
rect 6453 3299 6519 3302
rect 234797 3299 234863 3302
rect 295057 3362 295123 3365
rect 583385 3362 583451 3365
rect 295057 3360 583451 3362
rect 295057 3304 295062 3360
rect 295118 3304 583390 3360
rect 583446 3304 583451 3360
rect 295057 3302 583451 3304
rect 295057 3299 295123 3302
rect 583385 3299 583451 3302
<< via3 >>
rect 237236 377300 237300 377364
rect 238524 377300 238588 377364
rect 241284 377360 241348 377364
rect 241284 377304 241298 377360
rect 241298 377304 241348 377360
rect 241284 377300 241348 377304
rect 242756 377360 242820 377364
rect 242756 377304 242770 377360
rect 242770 377304 242820 377360
rect 242756 377300 242820 377304
rect 244044 377360 244108 377364
rect 244044 377304 244058 377360
rect 244058 377304 244108 377360
rect 244044 377300 244108 377304
rect 285812 377300 285876 377364
rect 287100 377300 287164 377364
rect 288388 377300 288452 377364
rect 290596 377300 290660 377364
rect 291148 377360 291212 377364
rect 291148 377304 291198 377360
rect 291198 377304 291212 377360
rect 291148 377300 291212 377304
rect 292620 377300 292684 377364
rect 285812 255172 285876 255236
rect 244044 218044 244108 218108
rect 287100 202812 287164 202876
rect 242756 178060 242820 178124
rect 290596 150316 290660 150380
rect 241284 138076 241348 138140
rect 288388 137940 288452 138004
rect 291148 97820 291212 97884
rect 238524 59332 238588 59396
rect 292620 59196 292684 59260
rect 237236 19348 237300 19412
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711002 -8694 711558
rect -8138 711002 -8106 711558
rect -8726 680614 -8106 711002
rect -8726 680058 -8694 680614
rect -8138 680058 -8106 680614
rect -8726 644614 -8106 680058
rect -8726 644058 -8694 644614
rect -8138 644058 -8106 644614
rect -8726 608614 -8106 644058
rect -8726 608058 -8694 608614
rect -8138 608058 -8106 608614
rect -8726 572614 -8106 608058
rect -8726 572058 -8694 572614
rect -8138 572058 -8106 572614
rect -8726 536614 -8106 572058
rect -8726 536058 -8694 536614
rect -8138 536058 -8106 536614
rect -8726 500614 -8106 536058
rect -8726 500058 -8694 500614
rect -8138 500058 -8106 500614
rect -8726 464614 -8106 500058
rect -8726 464058 -8694 464614
rect -8138 464058 -8106 464614
rect -8726 428614 -8106 464058
rect -8726 428058 -8694 428614
rect -8138 428058 -8106 428614
rect -8726 392614 -8106 428058
rect -8726 392058 -8694 392614
rect -8138 392058 -8106 392614
rect -8726 356614 -8106 392058
rect -8726 356058 -8694 356614
rect -8138 356058 -8106 356614
rect -8726 320614 -8106 356058
rect -8726 320058 -8694 320614
rect -8138 320058 -8106 320614
rect -8726 284614 -8106 320058
rect -8726 284058 -8694 284614
rect -8138 284058 -8106 284614
rect -8726 248614 -8106 284058
rect -8726 248058 -8694 248614
rect -8138 248058 -8106 248614
rect -8726 212614 -8106 248058
rect -8726 212058 -8694 212614
rect -8138 212058 -8106 212614
rect -8726 176614 -8106 212058
rect -8726 176058 -8694 176614
rect -8138 176058 -8106 176614
rect -8726 140614 -8106 176058
rect -8726 140058 -8694 140614
rect -8138 140058 -8106 140614
rect -8726 104614 -8106 140058
rect -8726 104058 -8694 104614
rect -8138 104058 -8106 104614
rect -8726 68614 -8106 104058
rect -8726 68058 -8694 68614
rect -8138 68058 -8106 68614
rect -8726 32614 -8106 68058
rect -8726 32058 -8694 32614
rect -8138 32058 -8106 32614
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710042 -7734 710598
rect -7178 710042 -7146 710598
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710042 12986 710598
rect 13542 710042 13574 710598
rect -7766 698058 -7734 698614
rect -7178 698058 -7146 698614
rect -7766 662614 -7146 698058
rect -7766 662058 -7734 662614
rect -7178 662058 -7146 662614
rect -7766 626614 -7146 662058
rect -7766 626058 -7734 626614
rect -7178 626058 -7146 626614
rect -7766 590614 -7146 626058
rect -7766 590058 -7734 590614
rect -7178 590058 -7146 590614
rect -7766 554614 -7146 590058
rect -7766 554058 -7734 554614
rect -7178 554058 -7146 554614
rect -7766 518614 -7146 554058
rect -7766 518058 -7734 518614
rect -7178 518058 -7146 518614
rect -7766 482614 -7146 518058
rect -7766 482058 -7734 482614
rect -7178 482058 -7146 482614
rect -7766 446614 -7146 482058
rect -7766 446058 -7734 446614
rect -7178 446058 -7146 446614
rect -7766 410614 -7146 446058
rect -7766 410058 -7734 410614
rect -7178 410058 -7146 410614
rect -7766 374614 -7146 410058
rect -7766 374058 -7734 374614
rect -7178 374058 -7146 374614
rect -7766 338614 -7146 374058
rect -7766 338058 -7734 338614
rect -7178 338058 -7146 338614
rect -7766 302614 -7146 338058
rect -7766 302058 -7734 302614
rect -7178 302058 -7146 302614
rect -7766 266614 -7146 302058
rect -7766 266058 -7734 266614
rect -7178 266058 -7146 266614
rect -7766 230614 -7146 266058
rect -7766 230058 -7734 230614
rect -7178 230058 -7146 230614
rect -7766 194614 -7146 230058
rect -7766 194058 -7734 194614
rect -7178 194058 -7146 194614
rect -7766 158614 -7146 194058
rect -7766 158058 -7734 158614
rect -7178 158058 -7146 158614
rect -7766 122614 -7146 158058
rect -7766 122058 -7734 122614
rect -7178 122058 -7146 122614
rect -7766 86614 -7146 122058
rect -7766 86058 -7734 86614
rect -7178 86058 -7146 86614
rect -7766 50614 -7146 86058
rect -7766 50058 -7734 50614
rect -7178 50058 -7146 50614
rect -7766 14614 -7146 50058
rect -7766 14058 -7734 14614
rect -7178 14058 -7146 14614
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709082 -6774 709638
rect -6218 709082 -6186 709638
rect -6806 676894 -6186 709082
rect -6806 676338 -6774 676894
rect -6218 676338 -6186 676894
rect -6806 640894 -6186 676338
rect -6806 640338 -6774 640894
rect -6218 640338 -6186 640894
rect -6806 604894 -6186 640338
rect -6806 604338 -6774 604894
rect -6218 604338 -6186 604894
rect -6806 568894 -6186 604338
rect -6806 568338 -6774 568894
rect -6218 568338 -6186 568894
rect -6806 532894 -6186 568338
rect -6806 532338 -6774 532894
rect -6218 532338 -6186 532894
rect -6806 496894 -6186 532338
rect -6806 496338 -6774 496894
rect -6218 496338 -6186 496894
rect -6806 460894 -6186 496338
rect -6806 460338 -6774 460894
rect -6218 460338 -6186 460894
rect -6806 424894 -6186 460338
rect -6806 424338 -6774 424894
rect -6218 424338 -6186 424894
rect -6806 388894 -6186 424338
rect -6806 388338 -6774 388894
rect -6218 388338 -6186 388894
rect -6806 352894 -6186 388338
rect -6806 352338 -6774 352894
rect -6218 352338 -6186 352894
rect -6806 316894 -6186 352338
rect -6806 316338 -6774 316894
rect -6218 316338 -6186 316894
rect -6806 280894 -6186 316338
rect -6806 280338 -6774 280894
rect -6218 280338 -6186 280894
rect -6806 244894 -6186 280338
rect -6806 244338 -6774 244894
rect -6218 244338 -6186 244894
rect -6806 208894 -6186 244338
rect -6806 208338 -6774 208894
rect -6218 208338 -6186 208894
rect -6806 172894 -6186 208338
rect -6806 172338 -6774 172894
rect -6218 172338 -6186 172894
rect -6806 136894 -6186 172338
rect -6806 136338 -6774 136894
rect -6218 136338 -6186 136894
rect -6806 100894 -6186 136338
rect -6806 100338 -6774 100894
rect -6218 100338 -6186 100894
rect -6806 64894 -6186 100338
rect -6806 64338 -6774 64894
rect -6218 64338 -6186 64894
rect -6806 28894 -6186 64338
rect -6806 28338 -6774 28894
rect -6218 28338 -6186 28894
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708122 -5814 708678
rect -5258 708122 -5226 708678
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708122 9266 708678
rect 9822 708122 9854 708678
rect -5846 694338 -5814 694894
rect -5258 694338 -5226 694894
rect -5846 658894 -5226 694338
rect -5846 658338 -5814 658894
rect -5258 658338 -5226 658894
rect -5846 622894 -5226 658338
rect -5846 622338 -5814 622894
rect -5258 622338 -5226 622894
rect -5846 586894 -5226 622338
rect -5846 586338 -5814 586894
rect -5258 586338 -5226 586894
rect -5846 550894 -5226 586338
rect -5846 550338 -5814 550894
rect -5258 550338 -5226 550894
rect -5846 514894 -5226 550338
rect -5846 514338 -5814 514894
rect -5258 514338 -5226 514894
rect -5846 478894 -5226 514338
rect -5846 478338 -5814 478894
rect -5258 478338 -5226 478894
rect -5846 442894 -5226 478338
rect -5846 442338 -5814 442894
rect -5258 442338 -5226 442894
rect -5846 406894 -5226 442338
rect -5846 406338 -5814 406894
rect -5258 406338 -5226 406894
rect -5846 370894 -5226 406338
rect -5846 370338 -5814 370894
rect -5258 370338 -5226 370894
rect -5846 334894 -5226 370338
rect -5846 334338 -5814 334894
rect -5258 334338 -5226 334894
rect -5846 298894 -5226 334338
rect -5846 298338 -5814 298894
rect -5258 298338 -5226 298894
rect -5846 262894 -5226 298338
rect -5846 262338 -5814 262894
rect -5258 262338 -5226 262894
rect -5846 226894 -5226 262338
rect -5846 226338 -5814 226894
rect -5258 226338 -5226 226894
rect -5846 190894 -5226 226338
rect -5846 190338 -5814 190894
rect -5258 190338 -5226 190894
rect -5846 154894 -5226 190338
rect -5846 154338 -5814 154894
rect -5258 154338 -5226 154894
rect -5846 118894 -5226 154338
rect -5846 118338 -5814 118894
rect -5258 118338 -5226 118894
rect -5846 82894 -5226 118338
rect -5846 82338 -5814 82894
rect -5258 82338 -5226 82894
rect -5846 46894 -5226 82338
rect -5846 46338 -5814 46894
rect -5258 46338 -5226 46894
rect -5846 10894 -5226 46338
rect -5846 10338 -5814 10894
rect -5258 10338 -5226 10894
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707162 -4854 707718
rect -4298 707162 -4266 707718
rect -4886 673174 -4266 707162
rect -4886 672618 -4854 673174
rect -4298 672618 -4266 673174
rect -4886 637174 -4266 672618
rect -4886 636618 -4854 637174
rect -4298 636618 -4266 637174
rect -4886 601174 -4266 636618
rect -4886 600618 -4854 601174
rect -4298 600618 -4266 601174
rect -4886 565174 -4266 600618
rect -4886 564618 -4854 565174
rect -4298 564618 -4266 565174
rect -4886 529174 -4266 564618
rect -4886 528618 -4854 529174
rect -4298 528618 -4266 529174
rect -4886 493174 -4266 528618
rect -4886 492618 -4854 493174
rect -4298 492618 -4266 493174
rect -4886 457174 -4266 492618
rect -4886 456618 -4854 457174
rect -4298 456618 -4266 457174
rect -4886 421174 -4266 456618
rect -4886 420618 -4854 421174
rect -4298 420618 -4266 421174
rect -4886 385174 -4266 420618
rect -4886 384618 -4854 385174
rect -4298 384618 -4266 385174
rect -4886 349174 -4266 384618
rect -4886 348618 -4854 349174
rect -4298 348618 -4266 349174
rect -4886 313174 -4266 348618
rect -4886 312618 -4854 313174
rect -4298 312618 -4266 313174
rect -4886 277174 -4266 312618
rect -4886 276618 -4854 277174
rect -4298 276618 -4266 277174
rect -4886 241174 -4266 276618
rect -4886 240618 -4854 241174
rect -4298 240618 -4266 241174
rect -4886 205174 -4266 240618
rect -4886 204618 -4854 205174
rect -4298 204618 -4266 205174
rect -4886 169174 -4266 204618
rect -4886 168618 -4854 169174
rect -4298 168618 -4266 169174
rect -4886 133174 -4266 168618
rect -4886 132618 -4854 133174
rect -4298 132618 -4266 133174
rect -4886 97174 -4266 132618
rect -4886 96618 -4854 97174
rect -4298 96618 -4266 97174
rect -4886 61174 -4266 96618
rect -4886 60618 -4854 61174
rect -4298 60618 -4266 61174
rect -4886 25174 -4266 60618
rect -4886 24618 -4854 25174
rect -4298 24618 -4266 25174
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706202 -3894 706758
rect -3338 706202 -3306 706758
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706202 5546 706758
rect 6102 706202 6134 706758
rect -3926 690618 -3894 691174
rect -3338 690618 -3306 691174
rect -3926 655174 -3306 690618
rect -3926 654618 -3894 655174
rect -3338 654618 -3306 655174
rect -3926 619174 -3306 654618
rect -3926 618618 -3894 619174
rect -3338 618618 -3306 619174
rect -3926 583174 -3306 618618
rect -3926 582618 -3894 583174
rect -3338 582618 -3306 583174
rect -3926 547174 -3306 582618
rect -3926 546618 -3894 547174
rect -3338 546618 -3306 547174
rect -3926 511174 -3306 546618
rect -3926 510618 -3894 511174
rect -3338 510618 -3306 511174
rect -3926 475174 -3306 510618
rect -3926 474618 -3894 475174
rect -3338 474618 -3306 475174
rect -3926 439174 -3306 474618
rect -3926 438618 -3894 439174
rect -3338 438618 -3306 439174
rect -3926 403174 -3306 438618
rect -3926 402618 -3894 403174
rect -3338 402618 -3306 403174
rect -3926 367174 -3306 402618
rect -3926 366618 -3894 367174
rect -3338 366618 -3306 367174
rect -3926 331174 -3306 366618
rect -3926 330618 -3894 331174
rect -3338 330618 -3306 331174
rect -3926 295174 -3306 330618
rect -3926 294618 -3894 295174
rect -3338 294618 -3306 295174
rect -3926 259174 -3306 294618
rect -3926 258618 -3894 259174
rect -3338 258618 -3306 259174
rect -3926 223174 -3306 258618
rect -3926 222618 -3894 223174
rect -3338 222618 -3306 223174
rect -3926 187174 -3306 222618
rect -3926 186618 -3894 187174
rect -3338 186618 -3306 187174
rect -3926 151174 -3306 186618
rect -3926 150618 -3894 151174
rect -3338 150618 -3306 151174
rect -3926 115174 -3306 150618
rect -3926 114618 -3894 115174
rect -3338 114618 -3306 115174
rect -3926 79174 -3306 114618
rect -3926 78618 -3894 79174
rect -3338 78618 -3306 79174
rect -3926 43174 -3306 78618
rect -3926 42618 -3894 43174
rect -3338 42618 -3306 43174
rect -3926 7174 -3306 42618
rect -3926 6618 -3894 7174
rect -3338 6618 -3306 7174
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705242 -2934 705798
rect -2378 705242 -2346 705798
rect -2966 669454 -2346 705242
rect -2966 668898 -2934 669454
rect -2378 668898 -2346 669454
rect -2966 633454 -2346 668898
rect -2966 632898 -2934 633454
rect -2378 632898 -2346 633454
rect -2966 597454 -2346 632898
rect -2966 596898 -2934 597454
rect -2378 596898 -2346 597454
rect -2966 561454 -2346 596898
rect -2966 560898 -2934 561454
rect -2378 560898 -2346 561454
rect -2966 525454 -2346 560898
rect -2966 524898 -2934 525454
rect -2378 524898 -2346 525454
rect -2966 489454 -2346 524898
rect -2966 488898 -2934 489454
rect -2378 488898 -2346 489454
rect -2966 453454 -2346 488898
rect -2966 452898 -2934 453454
rect -2378 452898 -2346 453454
rect -2966 417454 -2346 452898
rect -2966 416898 -2934 417454
rect -2378 416898 -2346 417454
rect -2966 381454 -2346 416898
rect -2966 380898 -2934 381454
rect -2378 380898 -2346 381454
rect -2966 345454 -2346 380898
rect -2966 344898 -2934 345454
rect -2378 344898 -2346 345454
rect -2966 309454 -2346 344898
rect -2966 308898 -2934 309454
rect -2378 308898 -2346 309454
rect -2966 273454 -2346 308898
rect -2966 272898 -2934 273454
rect -2378 272898 -2346 273454
rect -2966 237454 -2346 272898
rect -2966 236898 -2934 237454
rect -2378 236898 -2346 237454
rect -2966 201454 -2346 236898
rect -2966 200898 -2934 201454
rect -2378 200898 -2346 201454
rect -2966 165454 -2346 200898
rect -2966 164898 -2934 165454
rect -2378 164898 -2346 165454
rect -2966 129454 -2346 164898
rect -2966 128898 -2934 129454
rect -2378 128898 -2346 129454
rect -2966 93454 -2346 128898
rect -2966 92898 -2934 93454
rect -2378 92898 -2346 93454
rect -2966 57454 -2346 92898
rect -2966 56898 -2934 57454
rect -2378 56898 -2346 57454
rect -2966 21454 -2346 56898
rect -2966 20898 -2934 21454
rect -2378 20898 -2346 21454
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704282 -1974 704838
rect -1418 704282 -1386 704838
rect -2006 687454 -1386 704282
rect -2006 686898 -1974 687454
rect -1418 686898 -1386 687454
rect -2006 651454 -1386 686898
rect -2006 650898 -1974 651454
rect -1418 650898 -1386 651454
rect -2006 615454 -1386 650898
rect -2006 614898 -1974 615454
rect -1418 614898 -1386 615454
rect -2006 579454 -1386 614898
rect -2006 578898 -1974 579454
rect -1418 578898 -1386 579454
rect -2006 543454 -1386 578898
rect -2006 542898 -1974 543454
rect -1418 542898 -1386 543454
rect -2006 507454 -1386 542898
rect -2006 506898 -1974 507454
rect -1418 506898 -1386 507454
rect -2006 471454 -1386 506898
rect -2006 470898 -1974 471454
rect -1418 470898 -1386 471454
rect -2006 435454 -1386 470898
rect -2006 434898 -1974 435454
rect -1418 434898 -1386 435454
rect -2006 399454 -1386 434898
rect -2006 398898 -1974 399454
rect -1418 398898 -1386 399454
rect -2006 363454 -1386 398898
rect -2006 362898 -1974 363454
rect -1418 362898 -1386 363454
rect -2006 327454 -1386 362898
rect -2006 326898 -1974 327454
rect -1418 326898 -1386 327454
rect -2006 291454 -1386 326898
rect -2006 290898 -1974 291454
rect -1418 290898 -1386 291454
rect -2006 255454 -1386 290898
rect -2006 254898 -1974 255454
rect -1418 254898 -1386 255454
rect -2006 219454 -1386 254898
rect -2006 218898 -1974 219454
rect -1418 218898 -1386 219454
rect -2006 183454 -1386 218898
rect -2006 182898 -1974 183454
rect -1418 182898 -1386 183454
rect -2006 147454 -1386 182898
rect -2006 146898 -1974 147454
rect -1418 146898 -1386 147454
rect -2006 111454 -1386 146898
rect -2006 110898 -1974 111454
rect -1418 110898 -1386 111454
rect -2006 75454 -1386 110898
rect -2006 74898 -1974 75454
rect -1418 74898 -1386 75454
rect -2006 39454 -1386 74898
rect -2006 38898 -1974 39454
rect -1418 38898 -1386 39454
rect -2006 3454 -1386 38898
rect -2006 2898 -1974 3454
rect -1418 2898 -1386 3454
rect -2006 -346 -1386 2898
rect -2006 -902 -1974 -346
rect -1418 -902 -1386 -346
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704282 1826 704838
rect 2382 704282 2414 704838
rect 1794 687454 2414 704282
rect 1794 686898 1826 687454
rect 2382 686898 2414 687454
rect 1794 651454 2414 686898
rect 1794 650898 1826 651454
rect 2382 650898 2414 651454
rect 1794 615454 2414 650898
rect 1794 614898 1826 615454
rect 2382 614898 2414 615454
rect 1794 579454 2414 614898
rect 1794 578898 1826 579454
rect 2382 578898 2414 579454
rect 1794 543454 2414 578898
rect 1794 542898 1826 543454
rect 2382 542898 2414 543454
rect 1794 507454 2414 542898
rect 1794 506898 1826 507454
rect 2382 506898 2414 507454
rect 1794 471454 2414 506898
rect 1794 470898 1826 471454
rect 2382 470898 2414 471454
rect 1794 435454 2414 470898
rect 1794 434898 1826 435454
rect 2382 434898 2414 435454
rect 1794 399454 2414 434898
rect 1794 398898 1826 399454
rect 2382 398898 2414 399454
rect 1794 363454 2414 398898
rect 1794 362898 1826 363454
rect 2382 362898 2414 363454
rect 1794 327454 2414 362898
rect 1794 326898 1826 327454
rect 2382 326898 2414 327454
rect 1794 291454 2414 326898
rect 1794 290898 1826 291454
rect 2382 290898 2414 291454
rect 1794 255454 2414 290898
rect 1794 254898 1826 255454
rect 2382 254898 2414 255454
rect 1794 219454 2414 254898
rect 1794 218898 1826 219454
rect 2382 218898 2414 219454
rect 1794 183454 2414 218898
rect 1794 182898 1826 183454
rect 2382 182898 2414 183454
rect 1794 147454 2414 182898
rect 1794 146898 1826 147454
rect 2382 146898 2414 147454
rect 1794 111454 2414 146898
rect 1794 110898 1826 111454
rect 2382 110898 2414 111454
rect 1794 75454 2414 110898
rect 1794 74898 1826 75454
rect 2382 74898 2414 75454
rect 1794 39454 2414 74898
rect 1794 38898 1826 39454
rect 2382 38898 2414 39454
rect 1794 3454 2414 38898
rect 1794 2898 1826 3454
rect 2382 2898 2414 3454
rect 1794 -346 2414 2898
rect 1794 -902 1826 -346
rect 2382 -902 2414 -346
rect -2966 -1862 -2934 -1306
rect -2378 -1862 -2346 -1306
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690618 5546 691174
rect 6102 690618 6134 691174
rect 5514 655174 6134 690618
rect 5514 654618 5546 655174
rect 6102 654618 6134 655174
rect 5514 619174 6134 654618
rect 5514 618618 5546 619174
rect 6102 618618 6134 619174
rect 5514 583174 6134 618618
rect 5514 582618 5546 583174
rect 6102 582618 6134 583174
rect 5514 547174 6134 582618
rect 5514 546618 5546 547174
rect 6102 546618 6134 547174
rect 5514 511174 6134 546618
rect 5514 510618 5546 511174
rect 6102 510618 6134 511174
rect 5514 475174 6134 510618
rect 5514 474618 5546 475174
rect 6102 474618 6134 475174
rect 5514 439174 6134 474618
rect 5514 438618 5546 439174
rect 6102 438618 6134 439174
rect 5514 403174 6134 438618
rect 5514 402618 5546 403174
rect 6102 402618 6134 403174
rect 5514 367174 6134 402618
rect 5514 366618 5546 367174
rect 6102 366618 6134 367174
rect 5514 331174 6134 366618
rect 5514 330618 5546 331174
rect 6102 330618 6134 331174
rect 5514 295174 6134 330618
rect 5514 294618 5546 295174
rect 6102 294618 6134 295174
rect 5514 259174 6134 294618
rect 5514 258618 5546 259174
rect 6102 258618 6134 259174
rect 5514 223174 6134 258618
rect 5514 222618 5546 223174
rect 6102 222618 6134 223174
rect 5514 187174 6134 222618
rect 5514 186618 5546 187174
rect 6102 186618 6134 187174
rect 5514 151174 6134 186618
rect 5514 150618 5546 151174
rect 6102 150618 6134 151174
rect 5514 115174 6134 150618
rect 5514 114618 5546 115174
rect 6102 114618 6134 115174
rect 5514 79174 6134 114618
rect 5514 78618 5546 79174
rect 6102 78618 6134 79174
rect 5514 43174 6134 78618
rect 5514 42618 5546 43174
rect 6102 42618 6134 43174
rect 5514 7174 6134 42618
rect 5514 6618 5546 7174
rect 6102 6618 6134 7174
rect -3926 -2822 -3894 -2266
rect -3338 -2822 -3306 -2266
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2822 5546 -2266
rect 6102 -2822 6134 -2266
rect -4886 -3782 -4854 -3226
rect -4298 -3782 -4266 -3226
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694338 9266 694894
rect 9822 694338 9854 694894
rect 9234 658894 9854 694338
rect 9234 658338 9266 658894
rect 9822 658338 9854 658894
rect 9234 622894 9854 658338
rect 9234 622338 9266 622894
rect 9822 622338 9854 622894
rect 9234 586894 9854 622338
rect 9234 586338 9266 586894
rect 9822 586338 9854 586894
rect 9234 550894 9854 586338
rect 9234 550338 9266 550894
rect 9822 550338 9854 550894
rect 9234 514894 9854 550338
rect 9234 514338 9266 514894
rect 9822 514338 9854 514894
rect 9234 478894 9854 514338
rect 9234 478338 9266 478894
rect 9822 478338 9854 478894
rect 9234 442894 9854 478338
rect 9234 442338 9266 442894
rect 9822 442338 9854 442894
rect 9234 406894 9854 442338
rect 9234 406338 9266 406894
rect 9822 406338 9854 406894
rect 9234 370894 9854 406338
rect 9234 370338 9266 370894
rect 9822 370338 9854 370894
rect 9234 334894 9854 370338
rect 9234 334338 9266 334894
rect 9822 334338 9854 334894
rect 9234 298894 9854 334338
rect 9234 298338 9266 298894
rect 9822 298338 9854 298894
rect 9234 262894 9854 298338
rect 9234 262338 9266 262894
rect 9822 262338 9854 262894
rect 9234 226894 9854 262338
rect 9234 226338 9266 226894
rect 9822 226338 9854 226894
rect 9234 190894 9854 226338
rect 9234 190338 9266 190894
rect 9822 190338 9854 190894
rect 9234 154894 9854 190338
rect 9234 154338 9266 154894
rect 9822 154338 9854 154894
rect 9234 118894 9854 154338
rect 9234 118338 9266 118894
rect 9822 118338 9854 118894
rect 9234 82894 9854 118338
rect 9234 82338 9266 82894
rect 9822 82338 9854 82894
rect 9234 46894 9854 82338
rect 9234 46338 9266 46894
rect 9822 46338 9854 46894
rect 9234 10894 9854 46338
rect 9234 10338 9266 10894
rect 9822 10338 9854 10894
rect -5846 -4742 -5814 -4186
rect -5258 -4742 -5226 -4186
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4742 9266 -4186
rect 9822 -4742 9854 -4186
rect -6806 -5702 -6774 -5146
rect -6218 -5702 -6186 -5146
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711002 30986 711558
rect 31542 711002 31574 711558
rect 27234 709638 27854 709670
rect 27234 709082 27266 709638
rect 27822 709082 27854 709638
rect 23514 707718 24134 707750
rect 23514 707162 23546 707718
rect 24102 707162 24134 707718
rect 12954 698058 12986 698614
rect 13542 698058 13574 698614
rect 12954 662614 13574 698058
rect 12954 662058 12986 662614
rect 13542 662058 13574 662614
rect 12954 626614 13574 662058
rect 12954 626058 12986 626614
rect 13542 626058 13574 626614
rect 12954 590614 13574 626058
rect 12954 590058 12986 590614
rect 13542 590058 13574 590614
rect 12954 554614 13574 590058
rect 12954 554058 12986 554614
rect 13542 554058 13574 554614
rect 12954 518614 13574 554058
rect 12954 518058 12986 518614
rect 13542 518058 13574 518614
rect 12954 482614 13574 518058
rect 12954 482058 12986 482614
rect 13542 482058 13574 482614
rect 12954 446614 13574 482058
rect 12954 446058 12986 446614
rect 13542 446058 13574 446614
rect 12954 410614 13574 446058
rect 12954 410058 12986 410614
rect 13542 410058 13574 410614
rect 12954 374614 13574 410058
rect 12954 374058 12986 374614
rect 13542 374058 13574 374614
rect 12954 338614 13574 374058
rect 12954 338058 12986 338614
rect 13542 338058 13574 338614
rect 12954 302614 13574 338058
rect 12954 302058 12986 302614
rect 13542 302058 13574 302614
rect 12954 266614 13574 302058
rect 12954 266058 12986 266614
rect 13542 266058 13574 266614
rect 12954 230614 13574 266058
rect 12954 230058 12986 230614
rect 13542 230058 13574 230614
rect 12954 194614 13574 230058
rect 12954 194058 12986 194614
rect 13542 194058 13574 194614
rect 12954 158614 13574 194058
rect 12954 158058 12986 158614
rect 13542 158058 13574 158614
rect 12954 122614 13574 158058
rect 12954 122058 12986 122614
rect 13542 122058 13574 122614
rect 12954 86614 13574 122058
rect 12954 86058 12986 86614
rect 13542 86058 13574 86614
rect 12954 50614 13574 86058
rect 12954 50058 12986 50614
rect 13542 50058 13574 50614
rect 12954 14614 13574 50058
rect 12954 14058 12986 14614
rect 13542 14058 13574 14614
rect -7766 -6662 -7734 -6106
rect -7178 -6662 -7146 -6106
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705242 19826 705798
rect 20382 705242 20414 705798
rect 19794 669454 20414 705242
rect 19794 668898 19826 669454
rect 20382 668898 20414 669454
rect 19794 633454 20414 668898
rect 19794 632898 19826 633454
rect 20382 632898 20414 633454
rect 19794 597454 20414 632898
rect 19794 596898 19826 597454
rect 20382 596898 20414 597454
rect 19794 561454 20414 596898
rect 19794 560898 19826 561454
rect 20382 560898 20414 561454
rect 19794 525454 20414 560898
rect 19794 524898 19826 525454
rect 20382 524898 20414 525454
rect 19794 489454 20414 524898
rect 19794 488898 19826 489454
rect 20382 488898 20414 489454
rect 19794 453454 20414 488898
rect 19794 452898 19826 453454
rect 20382 452898 20414 453454
rect 19794 417454 20414 452898
rect 19794 416898 19826 417454
rect 20382 416898 20414 417454
rect 19794 381454 20414 416898
rect 19794 380898 19826 381454
rect 20382 380898 20414 381454
rect 19794 345454 20414 380898
rect 19794 344898 19826 345454
rect 20382 344898 20414 345454
rect 19794 309454 20414 344898
rect 19794 308898 19826 309454
rect 20382 308898 20414 309454
rect 19794 273454 20414 308898
rect 19794 272898 19826 273454
rect 20382 272898 20414 273454
rect 19794 237454 20414 272898
rect 19794 236898 19826 237454
rect 20382 236898 20414 237454
rect 19794 201454 20414 236898
rect 19794 200898 19826 201454
rect 20382 200898 20414 201454
rect 19794 165454 20414 200898
rect 19794 164898 19826 165454
rect 20382 164898 20414 165454
rect 19794 129454 20414 164898
rect 19794 128898 19826 129454
rect 20382 128898 20414 129454
rect 19794 93454 20414 128898
rect 19794 92898 19826 93454
rect 20382 92898 20414 93454
rect 19794 57454 20414 92898
rect 19794 56898 19826 57454
rect 20382 56898 20414 57454
rect 19794 21454 20414 56898
rect 19794 20898 19826 21454
rect 20382 20898 20414 21454
rect 19794 -1306 20414 20898
rect 19794 -1862 19826 -1306
rect 20382 -1862 20414 -1306
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672618 23546 673174
rect 24102 672618 24134 673174
rect 23514 637174 24134 672618
rect 23514 636618 23546 637174
rect 24102 636618 24134 637174
rect 23514 601174 24134 636618
rect 23514 600618 23546 601174
rect 24102 600618 24134 601174
rect 23514 565174 24134 600618
rect 23514 564618 23546 565174
rect 24102 564618 24134 565174
rect 23514 529174 24134 564618
rect 23514 528618 23546 529174
rect 24102 528618 24134 529174
rect 23514 493174 24134 528618
rect 23514 492618 23546 493174
rect 24102 492618 24134 493174
rect 23514 457174 24134 492618
rect 23514 456618 23546 457174
rect 24102 456618 24134 457174
rect 23514 421174 24134 456618
rect 23514 420618 23546 421174
rect 24102 420618 24134 421174
rect 23514 385174 24134 420618
rect 23514 384618 23546 385174
rect 24102 384618 24134 385174
rect 23514 349174 24134 384618
rect 23514 348618 23546 349174
rect 24102 348618 24134 349174
rect 23514 313174 24134 348618
rect 23514 312618 23546 313174
rect 24102 312618 24134 313174
rect 23514 277174 24134 312618
rect 23514 276618 23546 277174
rect 24102 276618 24134 277174
rect 23514 241174 24134 276618
rect 23514 240618 23546 241174
rect 24102 240618 24134 241174
rect 23514 205174 24134 240618
rect 23514 204618 23546 205174
rect 24102 204618 24134 205174
rect 23514 169174 24134 204618
rect 23514 168618 23546 169174
rect 24102 168618 24134 169174
rect 23514 133174 24134 168618
rect 23514 132618 23546 133174
rect 24102 132618 24134 133174
rect 23514 97174 24134 132618
rect 23514 96618 23546 97174
rect 24102 96618 24134 97174
rect 23514 61174 24134 96618
rect 23514 60618 23546 61174
rect 24102 60618 24134 61174
rect 23514 25174 24134 60618
rect 23514 24618 23546 25174
rect 24102 24618 24134 25174
rect 23514 -3226 24134 24618
rect 23514 -3782 23546 -3226
rect 24102 -3782 24134 -3226
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676338 27266 676894
rect 27822 676338 27854 676894
rect 27234 640894 27854 676338
rect 27234 640338 27266 640894
rect 27822 640338 27854 640894
rect 27234 604894 27854 640338
rect 27234 604338 27266 604894
rect 27822 604338 27854 604894
rect 27234 568894 27854 604338
rect 27234 568338 27266 568894
rect 27822 568338 27854 568894
rect 27234 532894 27854 568338
rect 27234 532338 27266 532894
rect 27822 532338 27854 532894
rect 27234 496894 27854 532338
rect 27234 496338 27266 496894
rect 27822 496338 27854 496894
rect 27234 460894 27854 496338
rect 27234 460338 27266 460894
rect 27822 460338 27854 460894
rect 27234 424894 27854 460338
rect 27234 424338 27266 424894
rect 27822 424338 27854 424894
rect 27234 388894 27854 424338
rect 27234 388338 27266 388894
rect 27822 388338 27854 388894
rect 27234 352894 27854 388338
rect 27234 352338 27266 352894
rect 27822 352338 27854 352894
rect 27234 316894 27854 352338
rect 27234 316338 27266 316894
rect 27822 316338 27854 316894
rect 27234 280894 27854 316338
rect 27234 280338 27266 280894
rect 27822 280338 27854 280894
rect 27234 244894 27854 280338
rect 27234 244338 27266 244894
rect 27822 244338 27854 244894
rect 27234 208894 27854 244338
rect 27234 208338 27266 208894
rect 27822 208338 27854 208894
rect 27234 172894 27854 208338
rect 27234 172338 27266 172894
rect 27822 172338 27854 172894
rect 27234 136894 27854 172338
rect 27234 136338 27266 136894
rect 27822 136338 27854 136894
rect 27234 100894 27854 136338
rect 27234 100338 27266 100894
rect 27822 100338 27854 100894
rect 27234 64894 27854 100338
rect 27234 64338 27266 64894
rect 27822 64338 27854 64894
rect 27234 28894 27854 64338
rect 27234 28338 27266 28894
rect 27822 28338 27854 28894
rect 27234 -5146 27854 28338
rect 27234 -5702 27266 -5146
rect 27822 -5702 27854 -5146
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710042 48986 710598
rect 49542 710042 49574 710598
rect 45234 708678 45854 709670
rect 45234 708122 45266 708678
rect 45822 708122 45854 708678
rect 41514 706758 42134 707750
rect 41514 706202 41546 706758
rect 42102 706202 42134 706758
rect 30954 680058 30986 680614
rect 31542 680058 31574 680614
rect 30954 644614 31574 680058
rect 30954 644058 30986 644614
rect 31542 644058 31574 644614
rect 30954 608614 31574 644058
rect 30954 608058 30986 608614
rect 31542 608058 31574 608614
rect 30954 572614 31574 608058
rect 30954 572058 30986 572614
rect 31542 572058 31574 572614
rect 30954 536614 31574 572058
rect 30954 536058 30986 536614
rect 31542 536058 31574 536614
rect 30954 500614 31574 536058
rect 30954 500058 30986 500614
rect 31542 500058 31574 500614
rect 30954 464614 31574 500058
rect 30954 464058 30986 464614
rect 31542 464058 31574 464614
rect 30954 428614 31574 464058
rect 30954 428058 30986 428614
rect 31542 428058 31574 428614
rect 30954 392614 31574 428058
rect 30954 392058 30986 392614
rect 31542 392058 31574 392614
rect 30954 356614 31574 392058
rect 30954 356058 30986 356614
rect 31542 356058 31574 356614
rect 30954 320614 31574 356058
rect 30954 320058 30986 320614
rect 31542 320058 31574 320614
rect 30954 284614 31574 320058
rect 30954 284058 30986 284614
rect 31542 284058 31574 284614
rect 30954 248614 31574 284058
rect 30954 248058 30986 248614
rect 31542 248058 31574 248614
rect 30954 212614 31574 248058
rect 30954 212058 30986 212614
rect 31542 212058 31574 212614
rect 30954 176614 31574 212058
rect 30954 176058 30986 176614
rect 31542 176058 31574 176614
rect 30954 140614 31574 176058
rect 30954 140058 30986 140614
rect 31542 140058 31574 140614
rect 30954 104614 31574 140058
rect 30954 104058 30986 104614
rect 31542 104058 31574 104614
rect 30954 68614 31574 104058
rect 30954 68058 30986 68614
rect 31542 68058 31574 68614
rect 30954 32614 31574 68058
rect 30954 32058 30986 32614
rect 31542 32058 31574 32614
rect 12954 -6662 12986 -6106
rect 13542 -6662 13574 -6106
rect -8726 -7622 -8694 -7066
rect -8138 -7622 -8106 -7066
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704282 37826 704838
rect 38382 704282 38414 704838
rect 37794 687454 38414 704282
rect 37794 686898 37826 687454
rect 38382 686898 38414 687454
rect 37794 651454 38414 686898
rect 37794 650898 37826 651454
rect 38382 650898 38414 651454
rect 37794 615454 38414 650898
rect 37794 614898 37826 615454
rect 38382 614898 38414 615454
rect 37794 579454 38414 614898
rect 37794 578898 37826 579454
rect 38382 578898 38414 579454
rect 37794 543454 38414 578898
rect 37794 542898 37826 543454
rect 38382 542898 38414 543454
rect 37794 507454 38414 542898
rect 37794 506898 37826 507454
rect 38382 506898 38414 507454
rect 37794 471454 38414 506898
rect 37794 470898 37826 471454
rect 38382 470898 38414 471454
rect 37794 435454 38414 470898
rect 37794 434898 37826 435454
rect 38382 434898 38414 435454
rect 37794 399454 38414 434898
rect 37794 398898 37826 399454
rect 38382 398898 38414 399454
rect 37794 363454 38414 398898
rect 37794 362898 37826 363454
rect 38382 362898 38414 363454
rect 37794 327454 38414 362898
rect 37794 326898 37826 327454
rect 38382 326898 38414 327454
rect 37794 291454 38414 326898
rect 37794 290898 37826 291454
rect 38382 290898 38414 291454
rect 37794 255454 38414 290898
rect 37794 254898 37826 255454
rect 38382 254898 38414 255454
rect 37794 219454 38414 254898
rect 37794 218898 37826 219454
rect 38382 218898 38414 219454
rect 37794 183454 38414 218898
rect 37794 182898 37826 183454
rect 38382 182898 38414 183454
rect 37794 147454 38414 182898
rect 37794 146898 37826 147454
rect 38382 146898 38414 147454
rect 37794 111454 38414 146898
rect 37794 110898 37826 111454
rect 38382 110898 38414 111454
rect 37794 75454 38414 110898
rect 37794 74898 37826 75454
rect 38382 74898 38414 75454
rect 37794 39454 38414 74898
rect 37794 38898 37826 39454
rect 38382 38898 38414 39454
rect 37794 3454 38414 38898
rect 37794 2898 37826 3454
rect 38382 2898 38414 3454
rect 37794 -346 38414 2898
rect 37794 -902 37826 -346
rect 38382 -902 38414 -346
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690618 41546 691174
rect 42102 690618 42134 691174
rect 41514 655174 42134 690618
rect 41514 654618 41546 655174
rect 42102 654618 42134 655174
rect 41514 619174 42134 654618
rect 41514 618618 41546 619174
rect 42102 618618 42134 619174
rect 41514 583174 42134 618618
rect 41514 582618 41546 583174
rect 42102 582618 42134 583174
rect 41514 547174 42134 582618
rect 41514 546618 41546 547174
rect 42102 546618 42134 547174
rect 41514 511174 42134 546618
rect 41514 510618 41546 511174
rect 42102 510618 42134 511174
rect 41514 475174 42134 510618
rect 41514 474618 41546 475174
rect 42102 474618 42134 475174
rect 41514 439174 42134 474618
rect 41514 438618 41546 439174
rect 42102 438618 42134 439174
rect 41514 403174 42134 438618
rect 41514 402618 41546 403174
rect 42102 402618 42134 403174
rect 41514 367174 42134 402618
rect 41514 366618 41546 367174
rect 42102 366618 42134 367174
rect 41514 331174 42134 366618
rect 41514 330618 41546 331174
rect 42102 330618 42134 331174
rect 41514 295174 42134 330618
rect 41514 294618 41546 295174
rect 42102 294618 42134 295174
rect 41514 259174 42134 294618
rect 41514 258618 41546 259174
rect 42102 258618 42134 259174
rect 41514 223174 42134 258618
rect 41514 222618 41546 223174
rect 42102 222618 42134 223174
rect 41514 187174 42134 222618
rect 41514 186618 41546 187174
rect 42102 186618 42134 187174
rect 41514 151174 42134 186618
rect 41514 150618 41546 151174
rect 42102 150618 42134 151174
rect 41514 115174 42134 150618
rect 41514 114618 41546 115174
rect 42102 114618 42134 115174
rect 41514 79174 42134 114618
rect 41514 78618 41546 79174
rect 42102 78618 42134 79174
rect 41514 43174 42134 78618
rect 41514 42618 41546 43174
rect 42102 42618 42134 43174
rect 41514 7174 42134 42618
rect 41514 6618 41546 7174
rect 42102 6618 42134 7174
rect 41514 -2266 42134 6618
rect 41514 -2822 41546 -2266
rect 42102 -2822 42134 -2266
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694338 45266 694894
rect 45822 694338 45854 694894
rect 45234 658894 45854 694338
rect 45234 658338 45266 658894
rect 45822 658338 45854 658894
rect 45234 622894 45854 658338
rect 45234 622338 45266 622894
rect 45822 622338 45854 622894
rect 45234 586894 45854 622338
rect 45234 586338 45266 586894
rect 45822 586338 45854 586894
rect 45234 550894 45854 586338
rect 45234 550338 45266 550894
rect 45822 550338 45854 550894
rect 45234 514894 45854 550338
rect 45234 514338 45266 514894
rect 45822 514338 45854 514894
rect 45234 478894 45854 514338
rect 45234 478338 45266 478894
rect 45822 478338 45854 478894
rect 45234 442894 45854 478338
rect 45234 442338 45266 442894
rect 45822 442338 45854 442894
rect 45234 406894 45854 442338
rect 45234 406338 45266 406894
rect 45822 406338 45854 406894
rect 45234 370894 45854 406338
rect 45234 370338 45266 370894
rect 45822 370338 45854 370894
rect 45234 334894 45854 370338
rect 45234 334338 45266 334894
rect 45822 334338 45854 334894
rect 45234 298894 45854 334338
rect 45234 298338 45266 298894
rect 45822 298338 45854 298894
rect 45234 262894 45854 298338
rect 45234 262338 45266 262894
rect 45822 262338 45854 262894
rect 45234 226894 45854 262338
rect 45234 226338 45266 226894
rect 45822 226338 45854 226894
rect 45234 190894 45854 226338
rect 45234 190338 45266 190894
rect 45822 190338 45854 190894
rect 45234 154894 45854 190338
rect 45234 154338 45266 154894
rect 45822 154338 45854 154894
rect 45234 118894 45854 154338
rect 45234 118338 45266 118894
rect 45822 118338 45854 118894
rect 45234 82894 45854 118338
rect 45234 82338 45266 82894
rect 45822 82338 45854 82894
rect 45234 46894 45854 82338
rect 45234 46338 45266 46894
rect 45822 46338 45854 46894
rect 45234 10894 45854 46338
rect 45234 10338 45266 10894
rect 45822 10338 45854 10894
rect 45234 -4186 45854 10338
rect 45234 -4742 45266 -4186
rect 45822 -4742 45854 -4186
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711002 66986 711558
rect 67542 711002 67574 711558
rect 63234 709638 63854 709670
rect 63234 709082 63266 709638
rect 63822 709082 63854 709638
rect 59514 707718 60134 707750
rect 59514 707162 59546 707718
rect 60102 707162 60134 707718
rect 48954 698058 48986 698614
rect 49542 698058 49574 698614
rect 48954 662614 49574 698058
rect 48954 662058 48986 662614
rect 49542 662058 49574 662614
rect 48954 626614 49574 662058
rect 48954 626058 48986 626614
rect 49542 626058 49574 626614
rect 48954 590614 49574 626058
rect 48954 590058 48986 590614
rect 49542 590058 49574 590614
rect 48954 554614 49574 590058
rect 48954 554058 48986 554614
rect 49542 554058 49574 554614
rect 48954 518614 49574 554058
rect 48954 518058 48986 518614
rect 49542 518058 49574 518614
rect 48954 482614 49574 518058
rect 48954 482058 48986 482614
rect 49542 482058 49574 482614
rect 48954 446614 49574 482058
rect 48954 446058 48986 446614
rect 49542 446058 49574 446614
rect 48954 410614 49574 446058
rect 48954 410058 48986 410614
rect 49542 410058 49574 410614
rect 48954 374614 49574 410058
rect 48954 374058 48986 374614
rect 49542 374058 49574 374614
rect 48954 338614 49574 374058
rect 48954 338058 48986 338614
rect 49542 338058 49574 338614
rect 48954 302614 49574 338058
rect 48954 302058 48986 302614
rect 49542 302058 49574 302614
rect 48954 266614 49574 302058
rect 48954 266058 48986 266614
rect 49542 266058 49574 266614
rect 48954 230614 49574 266058
rect 48954 230058 48986 230614
rect 49542 230058 49574 230614
rect 48954 194614 49574 230058
rect 48954 194058 48986 194614
rect 49542 194058 49574 194614
rect 48954 158614 49574 194058
rect 48954 158058 48986 158614
rect 49542 158058 49574 158614
rect 48954 122614 49574 158058
rect 48954 122058 48986 122614
rect 49542 122058 49574 122614
rect 48954 86614 49574 122058
rect 48954 86058 48986 86614
rect 49542 86058 49574 86614
rect 48954 50614 49574 86058
rect 48954 50058 48986 50614
rect 49542 50058 49574 50614
rect 48954 14614 49574 50058
rect 48954 14058 48986 14614
rect 49542 14058 49574 14614
rect 30954 -7622 30986 -7066
rect 31542 -7622 31574 -7066
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705242 55826 705798
rect 56382 705242 56414 705798
rect 55794 669454 56414 705242
rect 55794 668898 55826 669454
rect 56382 668898 56414 669454
rect 55794 633454 56414 668898
rect 55794 632898 55826 633454
rect 56382 632898 56414 633454
rect 55794 597454 56414 632898
rect 55794 596898 55826 597454
rect 56382 596898 56414 597454
rect 55794 561454 56414 596898
rect 55794 560898 55826 561454
rect 56382 560898 56414 561454
rect 55794 525454 56414 560898
rect 55794 524898 55826 525454
rect 56382 524898 56414 525454
rect 55794 489454 56414 524898
rect 55794 488898 55826 489454
rect 56382 488898 56414 489454
rect 55794 453454 56414 488898
rect 55794 452898 55826 453454
rect 56382 452898 56414 453454
rect 55794 417454 56414 452898
rect 55794 416898 55826 417454
rect 56382 416898 56414 417454
rect 55794 381454 56414 416898
rect 55794 380898 55826 381454
rect 56382 380898 56414 381454
rect 55794 345454 56414 380898
rect 55794 344898 55826 345454
rect 56382 344898 56414 345454
rect 55794 309454 56414 344898
rect 55794 308898 55826 309454
rect 56382 308898 56414 309454
rect 55794 273454 56414 308898
rect 55794 272898 55826 273454
rect 56382 272898 56414 273454
rect 55794 237454 56414 272898
rect 55794 236898 55826 237454
rect 56382 236898 56414 237454
rect 55794 201454 56414 236898
rect 55794 200898 55826 201454
rect 56382 200898 56414 201454
rect 55794 165454 56414 200898
rect 55794 164898 55826 165454
rect 56382 164898 56414 165454
rect 55794 129454 56414 164898
rect 55794 128898 55826 129454
rect 56382 128898 56414 129454
rect 55794 93454 56414 128898
rect 55794 92898 55826 93454
rect 56382 92898 56414 93454
rect 55794 57454 56414 92898
rect 55794 56898 55826 57454
rect 56382 56898 56414 57454
rect 55794 21454 56414 56898
rect 55794 20898 55826 21454
rect 56382 20898 56414 21454
rect 55794 -1306 56414 20898
rect 55794 -1862 55826 -1306
rect 56382 -1862 56414 -1306
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672618 59546 673174
rect 60102 672618 60134 673174
rect 59514 637174 60134 672618
rect 59514 636618 59546 637174
rect 60102 636618 60134 637174
rect 59514 601174 60134 636618
rect 59514 600618 59546 601174
rect 60102 600618 60134 601174
rect 59514 565174 60134 600618
rect 59514 564618 59546 565174
rect 60102 564618 60134 565174
rect 59514 529174 60134 564618
rect 59514 528618 59546 529174
rect 60102 528618 60134 529174
rect 59514 493174 60134 528618
rect 59514 492618 59546 493174
rect 60102 492618 60134 493174
rect 59514 457174 60134 492618
rect 59514 456618 59546 457174
rect 60102 456618 60134 457174
rect 59514 421174 60134 456618
rect 59514 420618 59546 421174
rect 60102 420618 60134 421174
rect 59514 385174 60134 420618
rect 59514 384618 59546 385174
rect 60102 384618 60134 385174
rect 59514 349174 60134 384618
rect 59514 348618 59546 349174
rect 60102 348618 60134 349174
rect 59514 313174 60134 348618
rect 59514 312618 59546 313174
rect 60102 312618 60134 313174
rect 59514 277174 60134 312618
rect 59514 276618 59546 277174
rect 60102 276618 60134 277174
rect 59514 241174 60134 276618
rect 59514 240618 59546 241174
rect 60102 240618 60134 241174
rect 59514 205174 60134 240618
rect 59514 204618 59546 205174
rect 60102 204618 60134 205174
rect 59514 169174 60134 204618
rect 59514 168618 59546 169174
rect 60102 168618 60134 169174
rect 59514 133174 60134 168618
rect 59514 132618 59546 133174
rect 60102 132618 60134 133174
rect 59514 97174 60134 132618
rect 59514 96618 59546 97174
rect 60102 96618 60134 97174
rect 59514 61174 60134 96618
rect 59514 60618 59546 61174
rect 60102 60618 60134 61174
rect 59514 25174 60134 60618
rect 59514 24618 59546 25174
rect 60102 24618 60134 25174
rect 59514 -3226 60134 24618
rect 59514 -3782 59546 -3226
rect 60102 -3782 60134 -3226
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676338 63266 676894
rect 63822 676338 63854 676894
rect 63234 640894 63854 676338
rect 63234 640338 63266 640894
rect 63822 640338 63854 640894
rect 63234 604894 63854 640338
rect 63234 604338 63266 604894
rect 63822 604338 63854 604894
rect 63234 568894 63854 604338
rect 63234 568338 63266 568894
rect 63822 568338 63854 568894
rect 63234 532894 63854 568338
rect 63234 532338 63266 532894
rect 63822 532338 63854 532894
rect 63234 496894 63854 532338
rect 63234 496338 63266 496894
rect 63822 496338 63854 496894
rect 63234 460894 63854 496338
rect 63234 460338 63266 460894
rect 63822 460338 63854 460894
rect 63234 424894 63854 460338
rect 63234 424338 63266 424894
rect 63822 424338 63854 424894
rect 63234 388894 63854 424338
rect 63234 388338 63266 388894
rect 63822 388338 63854 388894
rect 63234 352894 63854 388338
rect 63234 352338 63266 352894
rect 63822 352338 63854 352894
rect 63234 316894 63854 352338
rect 63234 316338 63266 316894
rect 63822 316338 63854 316894
rect 63234 280894 63854 316338
rect 63234 280338 63266 280894
rect 63822 280338 63854 280894
rect 63234 244894 63854 280338
rect 63234 244338 63266 244894
rect 63822 244338 63854 244894
rect 63234 208894 63854 244338
rect 63234 208338 63266 208894
rect 63822 208338 63854 208894
rect 63234 172894 63854 208338
rect 63234 172338 63266 172894
rect 63822 172338 63854 172894
rect 63234 136894 63854 172338
rect 63234 136338 63266 136894
rect 63822 136338 63854 136894
rect 63234 100894 63854 136338
rect 63234 100338 63266 100894
rect 63822 100338 63854 100894
rect 63234 64894 63854 100338
rect 63234 64338 63266 64894
rect 63822 64338 63854 64894
rect 63234 28894 63854 64338
rect 63234 28338 63266 28894
rect 63822 28338 63854 28894
rect 63234 -5146 63854 28338
rect 63234 -5702 63266 -5146
rect 63822 -5702 63854 -5146
rect 63234 -5734 63854 -5702
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710042 84986 710598
rect 85542 710042 85574 710598
rect 81234 708678 81854 709670
rect 81234 708122 81266 708678
rect 81822 708122 81854 708678
rect 77514 706758 78134 707750
rect 77514 706202 77546 706758
rect 78102 706202 78134 706758
rect 66954 680058 66986 680614
rect 67542 680058 67574 680614
rect 66954 644614 67574 680058
rect 66954 644058 66986 644614
rect 67542 644058 67574 644614
rect 66954 608614 67574 644058
rect 66954 608058 66986 608614
rect 67542 608058 67574 608614
rect 66954 572614 67574 608058
rect 66954 572058 66986 572614
rect 67542 572058 67574 572614
rect 66954 536614 67574 572058
rect 66954 536058 66986 536614
rect 67542 536058 67574 536614
rect 66954 500614 67574 536058
rect 66954 500058 66986 500614
rect 67542 500058 67574 500614
rect 66954 464614 67574 500058
rect 66954 464058 66986 464614
rect 67542 464058 67574 464614
rect 66954 428614 67574 464058
rect 66954 428058 66986 428614
rect 67542 428058 67574 428614
rect 66954 392614 67574 428058
rect 66954 392058 66986 392614
rect 67542 392058 67574 392614
rect 66954 356614 67574 392058
rect 66954 356058 66986 356614
rect 67542 356058 67574 356614
rect 66954 320614 67574 356058
rect 66954 320058 66986 320614
rect 67542 320058 67574 320614
rect 66954 284614 67574 320058
rect 66954 284058 66986 284614
rect 67542 284058 67574 284614
rect 66954 248614 67574 284058
rect 66954 248058 66986 248614
rect 67542 248058 67574 248614
rect 66954 212614 67574 248058
rect 66954 212058 66986 212614
rect 67542 212058 67574 212614
rect 66954 176614 67574 212058
rect 66954 176058 66986 176614
rect 67542 176058 67574 176614
rect 66954 140614 67574 176058
rect 66954 140058 66986 140614
rect 67542 140058 67574 140614
rect 66954 104614 67574 140058
rect 66954 104058 66986 104614
rect 67542 104058 67574 104614
rect 66954 68614 67574 104058
rect 66954 68058 66986 68614
rect 67542 68058 67574 68614
rect 66954 32614 67574 68058
rect 66954 32058 66986 32614
rect 67542 32058 67574 32614
rect 48954 -6662 48986 -6106
rect 49542 -6662 49574 -6106
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 704838 74414 705830
rect 73794 704282 73826 704838
rect 74382 704282 74414 704838
rect 73794 687454 74414 704282
rect 73794 686898 73826 687454
rect 74382 686898 74414 687454
rect 73794 651454 74414 686898
rect 73794 650898 73826 651454
rect 74382 650898 74414 651454
rect 73794 615454 74414 650898
rect 73794 614898 73826 615454
rect 74382 614898 74414 615454
rect 73794 579454 74414 614898
rect 73794 578898 73826 579454
rect 74382 578898 74414 579454
rect 73794 543454 74414 578898
rect 73794 542898 73826 543454
rect 74382 542898 74414 543454
rect 73794 507454 74414 542898
rect 73794 506898 73826 507454
rect 74382 506898 74414 507454
rect 73794 471454 74414 506898
rect 73794 470898 73826 471454
rect 74382 470898 74414 471454
rect 73794 435454 74414 470898
rect 73794 434898 73826 435454
rect 74382 434898 74414 435454
rect 73794 399454 74414 434898
rect 73794 398898 73826 399454
rect 74382 398898 74414 399454
rect 73794 363454 74414 398898
rect 73794 362898 73826 363454
rect 74382 362898 74414 363454
rect 73794 327454 74414 362898
rect 73794 326898 73826 327454
rect 74382 326898 74414 327454
rect 73794 291454 74414 326898
rect 73794 290898 73826 291454
rect 74382 290898 74414 291454
rect 73794 255454 74414 290898
rect 73794 254898 73826 255454
rect 74382 254898 74414 255454
rect 73794 219454 74414 254898
rect 73794 218898 73826 219454
rect 74382 218898 74414 219454
rect 73794 183454 74414 218898
rect 73794 182898 73826 183454
rect 74382 182898 74414 183454
rect 73794 147454 74414 182898
rect 73794 146898 73826 147454
rect 74382 146898 74414 147454
rect 73794 111454 74414 146898
rect 73794 110898 73826 111454
rect 74382 110898 74414 111454
rect 73794 75454 74414 110898
rect 73794 74898 73826 75454
rect 74382 74898 74414 75454
rect 73794 39454 74414 74898
rect 73794 38898 73826 39454
rect 74382 38898 74414 39454
rect 73794 3454 74414 38898
rect 73794 2898 73826 3454
rect 74382 2898 74414 3454
rect 73794 -346 74414 2898
rect 73794 -902 73826 -346
rect 74382 -902 74414 -346
rect 73794 -1894 74414 -902
rect 77514 691174 78134 706202
rect 77514 690618 77546 691174
rect 78102 690618 78134 691174
rect 77514 655174 78134 690618
rect 77514 654618 77546 655174
rect 78102 654618 78134 655174
rect 77514 619174 78134 654618
rect 77514 618618 77546 619174
rect 78102 618618 78134 619174
rect 77514 583174 78134 618618
rect 77514 582618 77546 583174
rect 78102 582618 78134 583174
rect 77514 547174 78134 582618
rect 77514 546618 77546 547174
rect 78102 546618 78134 547174
rect 77514 511174 78134 546618
rect 77514 510618 77546 511174
rect 78102 510618 78134 511174
rect 77514 475174 78134 510618
rect 77514 474618 77546 475174
rect 78102 474618 78134 475174
rect 77514 439174 78134 474618
rect 77514 438618 77546 439174
rect 78102 438618 78134 439174
rect 77514 403174 78134 438618
rect 77514 402618 77546 403174
rect 78102 402618 78134 403174
rect 77514 367174 78134 402618
rect 77514 366618 77546 367174
rect 78102 366618 78134 367174
rect 77514 331174 78134 366618
rect 77514 330618 77546 331174
rect 78102 330618 78134 331174
rect 77514 295174 78134 330618
rect 77514 294618 77546 295174
rect 78102 294618 78134 295174
rect 77514 259174 78134 294618
rect 77514 258618 77546 259174
rect 78102 258618 78134 259174
rect 77514 223174 78134 258618
rect 77514 222618 77546 223174
rect 78102 222618 78134 223174
rect 77514 187174 78134 222618
rect 77514 186618 77546 187174
rect 78102 186618 78134 187174
rect 77514 151174 78134 186618
rect 77514 150618 77546 151174
rect 78102 150618 78134 151174
rect 77514 115174 78134 150618
rect 77514 114618 77546 115174
rect 78102 114618 78134 115174
rect 77514 79174 78134 114618
rect 77514 78618 77546 79174
rect 78102 78618 78134 79174
rect 77514 43174 78134 78618
rect 77514 42618 77546 43174
rect 78102 42618 78134 43174
rect 77514 7174 78134 42618
rect 77514 6618 77546 7174
rect 78102 6618 78134 7174
rect 77514 -2266 78134 6618
rect 77514 -2822 77546 -2266
rect 78102 -2822 78134 -2266
rect 77514 -3814 78134 -2822
rect 81234 694894 81854 708122
rect 81234 694338 81266 694894
rect 81822 694338 81854 694894
rect 81234 658894 81854 694338
rect 81234 658338 81266 658894
rect 81822 658338 81854 658894
rect 81234 622894 81854 658338
rect 81234 622338 81266 622894
rect 81822 622338 81854 622894
rect 81234 586894 81854 622338
rect 81234 586338 81266 586894
rect 81822 586338 81854 586894
rect 81234 550894 81854 586338
rect 81234 550338 81266 550894
rect 81822 550338 81854 550894
rect 81234 514894 81854 550338
rect 81234 514338 81266 514894
rect 81822 514338 81854 514894
rect 81234 478894 81854 514338
rect 81234 478338 81266 478894
rect 81822 478338 81854 478894
rect 81234 442894 81854 478338
rect 81234 442338 81266 442894
rect 81822 442338 81854 442894
rect 81234 406894 81854 442338
rect 81234 406338 81266 406894
rect 81822 406338 81854 406894
rect 81234 370894 81854 406338
rect 81234 370338 81266 370894
rect 81822 370338 81854 370894
rect 81234 334894 81854 370338
rect 81234 334338 81266 334894
rect 81822 334338 81854 334894
rect 81234 298894 81854 334338
rect 81234 298338 81266 298894
rect 81822 298338 81854 298894
rect 81234 262894 81854 298338
rect 81234 262338 81266 262894
rect 81822 262338 81854 262894
rect 81234 226894 81854 262338
rect 81234 226338 81266 226894
rect 81822 226338 81854 226894
rect 81234 190894 81854 226338
rect 81234 190338 81266 190894
rect 81822 190338 81854 190894
rect 81234 154894 81854 190338
rect 81234 154338 81266 154894
rect 81822 154338 81854 154894
rect 81234 118894 81854 154338
rect 81234 118338 81266 118894
rect 81822 118338 81854 118894
rect 81234 82894 81854 118338
rect 81234 82338 81266 82894
rect 81822 82338 81854 82894
rect 81234 46894 81854 82338
rect 81234 46338 81266 46894
rect 81822 46338 81854 46894
rect 81234 10894 81854 46338
rect 81234 10338 81266 10894
rect 81822 10338 81854 10894
rect 81234 -4186 81854 10338
rect 81234 -4742 81266 -4186
rect 81822 -4742 81854 -4186
rect 81234 -5734 81854 -4742
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711002 102986 711558
rect 103542 711002 103574 711558
rect 99234 709638 99854 709670
rect 99234 709082 99266 709638
rect 99822 709082 99854 709638
rect 95514 707718 96134 707750
rect 95514 707162 95546 707718
rect 96102 707162 96134 707718
rect 84954 698058 84986 698614
rect 85542 698058 85574 698614
rect 84954 662614 85574 698058
rect 84954 662058 84986 662614
rect 85542 662058 85574 662614
rect 84954 626614 85574 662058
rect 84954 626058 84986 626614
rect 85542 626058 85574 626614
rect 84954 590614 85574 626058
rect 84954 590058 84986 590614
rect 85542 590058 85574 590614
rect 84954 554614 85574 590058
rect 84954 554058 84986 554614
rect 85542 554058 85574 554614
rect 84954 518614 85574 554058
rect 84954 518058 84986 518614
rect 85542 518058 85574 518614
rect 84954 482614 85574 518058
rect 84954 482058 84986 482614
rect 85542 482058 85574 482614
rect 84954 446614 85574 482058
rect 84954 446058 84986 446614
rect 85542 446058 85574 446614
rect 84954 410614 85574 446058
rect 84954 410058 84986 410614
rect 85542 410058 85574 410614
rect 84954 374614 85574 410058
rect 84954 374058 84986 374614
rect 85542 374058 85574 374614
rect 84954 338614 85574 374058
rect 84954 338058 84986 338614
rect 85542 338058 85574 338614
rect 84954 302614 85574 338058
rect 84954 302058 84986 302614
rect 85542 302058 85574 302614
rect 84954 266614 85574 302058
rect 84954 266058 84986 266614
rect 85542 266058 85574 266614
rect 84954 230614 85574 266058
rect 84954 230058 84986 230614
rect 85542 230058 85574 230614
rect 84954 194614 85574 230058
rect 84954 194058 84986 194614
rect 85542 194058 85574 194614
rect 84954 158614 85574 194058
rect 84954 158058 84986 158614
rect 85542 158058 85574 158614
rect 84954 122614 85574 158058
rect 84954 122058 84986 122614
rect 85542 122058 85574 122614
rect 84954 86614 85574 122058
rect 84954 86058 84986 86614
rect 85542 86058 85574 86614
rect 84954 50614 85574 86058
rect 84954 50058 84986 50614
rect 85542 50058 85574 50614
rect 84954 14614 85574 50058
rect 84954 14058 84986 14614
rect 85542 14058 85574 14614
rect 66954 -7622 66986 -7066
rect 67542 -7622 67574 -7066
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 705798 92414 705830
rect 91794 705242 91826 705798
rect 92382 705242 92414 705798
rect 91794 669454 92414 705242
rect 91794 668898 91826 669454
rect 92382 668898 92414 669454
rect 91794 633454 92414 668898
rect 91794 632898 91826 633454
rect 92382 632898 92414 633454
rect 91794 597454 92414 632898
rect 91794 596898 91826 597454
rect 92382 596898 92414 597454
rect 91794 561454 92414 596898
rect 91794 560898 91826 561454
rect 92382 560898 92414 561454
rect 91794 525454 92414 560898
rect 91794 524898 91826 525454
rect 92382 524898 92414 525454
rect 91794 489454 92414 524898
rect 91794 488898 91826 489454
rect 92382 488898 92414 489454
rect 91794 453454 92414 488898
rect 91794 452898 91826 453454
rect 92382 452898 92414 453454
rect 91794 417454 92414 452898
rect 91794 416898 91826 417454
rect 92382 416898 92414 417454
rect 91794 381454 92414 416898
rect 91794 380898 91826 381454
rect 92382 380898 92414 381454
rect 91794 345454 92414 380898
rect 91794 344898 91826 345454
rect 92382 344898 92414 345454
rect 91794 309454 92414 344898
rect 91794 308898 91826 309454
rect 92382 308898 92414 309454
rect 91794 273454 92414 308898
rect 91794 272898 91826 273454
rect 92382 272898 92414 273454
rect 91794 237454 92414 272898
rect 91794 236898 91826 237454
rect 92382 236898 92414 237454
rect 91794 201454 92414 236898
rect 91794 200898 91826 201454
rect 92382 200898 92414 201454
rect 91794 165454 92414 200898
rect 91794 164898 91826 165454
rect 92382 164898 92414 165454
rect 91794 129454 92414 164898
rect 91794 128898 91826 129454
rect 92382 128898 92414 129454
rect 91794 93454 92414 128898
rect 91794 92898 91826 93454
rect 92382 92898 92414 93454
rect 91794 57454 92414 92898
rect 91794 56898 91826 57454
rect 92382 56898 92414 57454
rect 91794 21454 92414 56898
rect 91794 20898 91826 21454
rect 92382 20898 92414 21454
rect 91794 -1306 92414 20898
rect 91794 -1862 91826 -1306
rect 92382 -1862 92414 -1306
rect 91794 -1894 92414 -1862
rect 95514 673174 96134 707162
rect 95514 672618 95546 673174
rect 96102 672618 96134 673174
rect 95514 637174 96134 672618
rect 95514 636618 95546 637174
rect 96102 636618 96134 637174
rect 95514 601174 96134 636618
rect 95514 600618 95546 601174
rect 96102 600618 96134 601174
rect 95514 565174 96134 600618
rect 95514 564618 95546 565174
rect 96102 564618 96134 565174
rect 95514 529174 96134 564618
rect 95514 528618 95546 529174
rect 96102 528618 96134 529174
rect 95514 493174 96134 528618
rect 95514 492618 95546 493174
rect 96102 492618 96134 493174
rect 95514 457174 96134 492618
rect 95514 456618 95546 457174
rect 96102 456618 96134 457174
rect 95514 421174 96134 456618
rect 95514 420618 95546 421174
rect 96102 420618 96134 421174
rect 95514 385174 96134 420618
rect 95514 384618 95546 385174
rect 96102 384618 96134 385174
rect 95514 349174 96134 384618
rect 95514 348618 95546 349174
rect 96102 348618 96134 349174
rect 95514 313174 96134 348618
rect 95514 312618 95546 313174
rect 96102 312618 96134 313174
rect 95514 277174 96134 312618
rect 95514 276618 95546 277174
rect 96102 276618 96134 277174
rect 95514 241174 96134 276618
rect 95514 240618 95546 241174
rect 96102 240618 96134 241174
rect 95514 205174 96134 240618
rect 95514 204618 95546 205174
rect 96102 204618 96134 205174
rect 95514 169174 96134 204618
rect 95514 168618 95546 169174
rect 96102 168618 96134 169174
rect 95514 133174 96134 168618
rect 95514 132618 95546 133174
rect 96102 132618 96134 133174
rect 95514 97174 96134 132618
rect 95514 96618 95546 97174
rect 96102 96618 96134 97174
rect 95514 61174 96134 96618
rect 95514 60618 95546 61174
rect 96102 60618 96134 61174
rect 95514 25174 96134 60618
rect 95514 24618 95546 25174
rect 96102 24618 96134 25174
rect 95514 -3226 96134 24618
rect 95514 -3782 95546 -3226
rect 96102 -3782 96134 -3226
rect 95514 -3814 96134 -3782
rect 99234 676894 99854 709082
rect 99234 676338 99266 676894
rect 99822 676338 99854 676894
rect 99234 640894 99854 676338
rect 99234 640338 99266 640894
rect 99822 640338 99854 640894
rect 99234 604894 99854 640338
rect 99234 604338 99266 604894
rect 99822 604338 99854 604894
rect 99234 568894 99854 604338
rect 99234 568338 99266 568894
rect 99822 568338 99854 568894
rect 99234 532894 99854 568338
rect 99234 532338 99266 532894
rect 99822 532338 99854 532894
rect 99234 496894 99854 532338
rect 99234 496338 99266 496894
rect 99822 496338 99854 496894
rect 99234 460894 99854 496338
rect 99234 460338 99266 460894
rect 99822 460338 99854 460894
rect 99234 424894 99854 460338
rect 99234 424338 99266 424894
rect 99822 424338 99854 424894
rect 99234 388894 99854 424338
rect 99234 388338 99266 388894
rect 99822 388338 99854 388894
rect 99234 352894 99854 388338
rect 99234 352338 99266 352894
rect 99822 352338 99854 352894
rect 99234 316894 99854 352338
rect 99234 316338 99266 316894
rect 99822 316338 99854 316894
rect 99234 280894 99854 316338
rect 99234 280338 99266 280894
rect 99822 280338 99854 280894
rect 99234 244894 99854 280338
rect 99234 244338 99266 244894
rect 99822 244338 99854 244894
rect 99234 208894 99854 244338
rect 99234 208338 99266 208894
rect 99822 208338 99854 208894
rect 99234 172894 99854 208338
rect 99234 172338 99266 172894
rect 99822 172338 99854 172894
rect 99234 136894 99854 172338
rect 99234 136338 99266 136894
rect 99822 136338 99854 136894
rect 99234 100894 99854 136338
rect 99234 100338 99266 100894
rect 99822 100338 99854 100894
rect 99234 64894 99854 100338
rect 99234 64338 99266 64894
rect 99822 64338 99854 64894
rect 99234 28894 99854 64338
rect 99234 28338 99266 28894
rect 99822 28338 99854 28894
rect 99234 -5146 99854 28338
rect 99234 -5702 99266 -5146
rect 99822 -5702 99854 -5146
rect 99234 -5734 99854 -5702
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710042 120986 710598
rect 121542 710042 121574 710598
rect 117234 708678 117854 709670
rect 117234 708122 117266 708678
rect 117822 708122 117854 708678
rect 113514 706758 114134 707750
rect 113514 706202 113546 706758
rect 114102 706202 114134 706758
rect 102954 680058 102986 680614
rect 103542 680058 103574 680614
rect 102954 644614 103574 680058
rect 102954 644058 102986 644614
rect 103542 644058 103574 644614
rect 102954 608614 103574 644058
rect 102954 608058 102986 608614
rect 103542 608058 103574 608614
rect 102954 572614 103574 608058
rect 102954 572058 102986 572614
rect 103542 572058 103574 572614
rect 102954 536614 103574 572058
rect 102954 536058 102986 536614
rect 103542 536058 103574 536614
rect 102954 500614 103574 536058
rect 102954 500058 102986 500614
rect 103542 500058 103574 500614
rect 102954 464614 103574 500058
rect 102954 464058 102986 464614
rect 103542 464058 103574 464614
rect 102954 428614 103574 464058
rect 102954 428058 102986 428614
rect 103542 428058 103574 428614
rect 102954 392614 103574 428058
rect 102954 392058 102986 392614
rect 103542 392058 103574 392614
rect 102954 356614 103574 392058
rect 102954 356058 102986 356614
rect 103542 356058 103574 356614
rect 102954 320614 103574 356058
rect 102954 320058 102986 320614
rect 103542 320058 103574 320614
rect 102954 284614 103574 320058
rect 102954 284058 102986 284614
rect 103542 284058 103574 284614
rect 102954 248614 103574 284058
rect 102954 248058 102986 248614
rect 103542 248058 103574 248614
rect 102954 212614 103574 248058
rect 102954 212058 102986 212614
rect 103542 212058 103574 212614
rect 102954 176614 103574 212058
rect 102954 176058 102986 176614
rect 103542 176058 103574 176614
rect 102954 140614 103574 176058
rect 102954 140058 102986 140614
rect 103542 140058 103574 140614
rect 102954 104614 103574 140058
rect 102954 104058 102986 104614
rect 103542 104058 103574 104614
rect 102954 68614 103574 104058
rect 102954 68058 102986 68614
rect 103542 68058 103574 68614
rect 102954 32614 103574 68058
rect 102954 32058 102986 32614
rect 103542 32058 103574 32614
rect 84954 -6662 84986 -6106
rect 85542 -6662 85574 -6106
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 704838 110414 705830
rect 109794 704282 109826 704838
rect 110382 704282 110414 704838
rect 109794 687454 110414 704282
rect 109794 686898 109826 687454
rect 110382 686898 110414 687454
rect 109794 651454 110414 686898
rect 109794 650898 109826 651454
rect 110382 650898 110414 651454
rect 109794 615454 110414 650898
rect 109794 614898 109826 615454
rect 110382 614898 110414 615454
rect 109794 579454 110414 614898
rect 109794 578898 109826 579454
rect 110382 578898 110414 579454
rect 109794 543454 110414 578898
rect 109794 542898 109826 543454
rect 110382 542898 110414 543454
rect 109794 507454 110414 542898
rect 109794 506898 109826 507454
rect 110382 506898 110414 507454
rect 109794 471454 110414 506898
rect 109794 470898 109826 471454
rect 110382 470898 110414 471454
rect 109794 435454 110414 470898
rect 109794 434898 109826 435454
rect 110382 434898 110414 435454
rect 109794 399454 110414 434898
rect 109794 398898 109826 399454
rect 110382 398898 110414 399454
rect 109794 363454 110414 398898
rect 109794 362898 109826 363454
rect 110382 362898 110414 363454
rect 109794 327454 110414 362898
rect 109794 326898 109826 327454
rect 110382 326898 110414 327454
rect 109794 291454 110414 326898
rect 109794 290898 109826 291454
rect 110382 290898 110414 291454
rect 109794 255454 110414 290898
rect 109794 254898 109826 255454
rect 110382 254898 110414 255454
rect 109794 219454 110414 254898
rect 109794 218898 109826 219454
rect 110382 218898 110414 219454
rect 109794 183454 110414 218898
rect 109794 182898 109826 183454
rect 110382 182898 110414 183454
rect 109794 147454 110414 182898
rect 109794 146898 109826 147454
rect 110382 146898 110414 147454
rect 109794 111454 110414 146898
rect 109794 110898 109826 111454
rect 110382 110898 110414 111454
rect 109794 75454 110414 110898
rect 109794 74898 109826 75454
rect 110382 74898 110414 75454
rect 109794 39454 110414 74898
rect 109794 38898 109826 39454
rect 110382 38898 110414 39454
rect 109794 3454 110414 38898
rect 109794 2898 109826 3454
rect 110382 2898 110414 3454
rect 109794 -346 110414 2898
rect 109794 -902 109826 -346
rect 110382 -902 110414 -346
rect 109794 -1894 110414 -902
rect 113514 691174 114134 706202
rect 113514 690618 113546 691174
rect 114102 690618 114134 691174
rect 113514 655174 114134 690618
rect 113514 654618 113546 655174
rect 114102 654618 114134 655174
rect 113514 619174 114134 654618
rect 113514 618618 113546 619174
rect 114102 618618 114134 619174
rect 113514 583174 114134 618618
rect 113514 582618 113546 583174
rect 114102 582618 114134 583174
rect 113514 547174 114134 582618
rect 113514 546618 113546 547174
rect 114102 546618 114134 547174
rect 113514 511174 114134 546618
rect 113514 510618 113546 511174
rect 114102 510618 114134 511174
rect 113514 475174 114134 510618
rect 113514 474618 113546 475174
rect 114102 474618 114134 475174
rect 113514 439174 114134 474618
rect 113514 438618 113546 439174
rect 114102 438618 114134 439174
rect 113514 403174 114134 438618
rect 113514 402618 113546 403174
rect 114102 402618 114134 403174
rect 113514 367174 114134 402618
rect 113514 366618 113546 367174
rect 114102 366618 114134 367174
rect 113514 331174 114134 366618
rect 113514 330618 113546 331174
rect 114102 330618 114134 331174
rect 113514 295174 114134 330618
rect 113514 294618 113546 295174
rect 114102 294618 114134 295174
rect 113514 259174 114134 294618
rect 113514 258618 113546 259174
rect 114102 258618 114134 259174
rect 113514 223174 114134 258618
rect 113514 222618 113546 223174
rect 114102 222618 114134 223174
rect 113514 187174 114134 222618
rect 113514 186618 113546 187174
rect 114102 186618 114134 187174
rect 113514 151174 114134 186618
rect 113514 150618 113546 151174
rect 114102 150618 114134 151174
rect 113514 115174 114134 150618
rect 113514 114618 113546 115174
rect 114102 114618 114134 115174
rect 113514 79174 114134 114618
rect 113514 78618 113546 79174
rect 114102 78618 114134 79174
rect 113514 43174 114134 78618
rect 113514 42618 113546 43174
rect 114102 42618 114134 43174
rect 113514 7174 114134 42618
rect 113514 6618 113546 7174
rect 114102 6618 114134 7174
rect 113514 -2266 114134 6618
rect 113514 -2822 113546 -2266
rect 114102 -2822 114134 -2266
rect 113514 -3814 114134 -2822
rect 117234 694894 117854 708122
rect 117234 694338 117266 694894
rect 117822 694338 117854 694894
rect 117234 658894 117854 694338
rect 117234 658338 117266 658894
rect 117822 658338 117854 658894
rect 117234 622894 117854 658338
rect 117234 622338 117266 622894
rect 117822 622338 117854 622894
rect 117234 586894 117854 622338
rect 117234 586338 117266 586894
rect 117822 586338 117854 586894
rect 117234 550894 117854 586338
rect 117234 550338 117266 550894
rect 117822 550338 117854 550894
rect 117234 514894 117854 550338
rect 117234 514338 117266 514894
rect 117822 514338 117854 514894
rect 117234 478894 117854 514338
rect 117234 478338 117266 478894
rect 117822 478338 117854 478894
rect 117234 442894 117854 478338
rect 117234 442338 117266 442894
rect 117822 442338 117854 442894
rect 117234 406894 117854 442338
rect 117234 406338 117266 406894
rect 117822 406338 117854 406894
rect 117234 370894 117854 406338
rect 117234 370338 117266 370894
rect 117822 370338 117854 370894
rect 117234 334894 117854 370338
rect 117234 334338 117266 334894
rect 117822 334338 117854 334894
rect 117234 298894 117854 334338
rect 117234 298338 117266 298894
rect 117822 298338 117854 298894
rect 117234 262894 117854 298338
rect 117234 262338 117266 262894
rect 117822 262338 117854 262894
rect 117234 226894 117854 262338
rect 117234 226338 117266 226894
rect 117822 226338 117854 226894
rect 117234 190894 117854 226338
rect 117234 190338 117266 190894
rect 117822 190338 117854 190894
rect 117234 154894 117854 190338
rect 117234 154338 117266 154894
rect 117822 154338 117854 154894
rect 117234 118894 117854 154338
rect 117234 118338 117266 118894
rect 117822 118338 117854 118894
rect 117234 82894 117854 118338
rect 117234 82338 117266 82894
rect 117822 82338 117854 82894
rect 117234 46894 117854 82338
rect 117234 46338 117266 46894
rect 117822 46338 117854 46894
rect 117234 10894 117854 46338
rect 117234 10338 117266 10894
rect 117822 10338 117854 10894
rect 117234 -4186 117854 10338
rect 117234 -4742 117266 -4186
rect 117822 -4742 117854 -4186
rect 117234 -5734 117854 -4742
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711002 138986 711558
rect 139542 711002 139574 711558
rect 135234 709638 135854 709670
rect 135234 709082 135266 709638
rect 135822 709082 135854 709638
rect 131514 707718 132134 707750
rect 131514 707162 131546 707718
rect 132102 707162 132134 707718
rect 120954 698058 120986 698614
rect 121542 698058 121574 698614
rect 120954 662614 121574 698058
rect 120954 662058 120986 662614
rect 121542 662058 121574 662614
rect 120954 626614 121574 662058
rect 120954 626058 120986 626614
rect 121542 626058 121574 626614
rect 120954 590614 121574 626058
rect 120954 590058 120986 590614
rect 121542 590058 121574 590614
rect 120954 554614 121574 590058
rect 120954 554058 120986 554614
rect 121542 554058 121574 554614
rect 120954 518614 121574 554058
rect 120954 518058 120986 518614
rect 121542 518058 121574 518614
rect 120954 482614 121574 518058
rect 120954 482058 120986 482614
rect 121542 482058 121574 482614
rect 120954 446614 121574 482058
rect 120954 446058 120986 446614
rect 121542 446058 121574 446614
rect 120954 410614 121574 446058
rect 120954 410058 120986 410614
rect 121542 410058 121574 410614
rect 120954 374614 121574 410058
rect 120954 374058 120986 374614
rect 121542 374058 121574 374614
rect 120954 338614 121574 374058
rect 120954 338058 120986 338614
rect 121542 338058 121574 338614
rect 120954 302614 121574 338058
rect 120954 302058 120986 302614
rect 121542 302058 121574 302614
rect 120954 266614 121574 302058
rect 120954 266058 120986 266614
rect 121542 266058 121574 266614
rect 120954 230614 121574 266058
rect 120954 230058 120986 230614
rect 121542 230058 121574 230614
rect 120954 194614 121574 230058
rect 120954 194058 120986 194614
rect 121542 194058 121574 194614
rect 120954 158614 121574 194058
rect 120954 158058 120986 158614
rect 121542 158058 121574 158614
rect 120954 122614 121574 158058
rect 120954 122058 120986 122614
rect 121542 122058 121574 122614
rect 120954 86614 121574 122058
rect 120954 86058 120986 86614
rect 121542 86058 121574 86614
rect 120954 50614 121574 86058
rect 120954 50058 120986 50614
rect 121542 50058 121574 50614
rect 120954 14614 121574 50058
rect 120954 14058 120986 14614
rect 121542 14058 121574 14614
rect 102954 -7622 102986 -7066
rect 103542 -7622 103574 -7066
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 705798 128414 705830
rect 127794 705242 127826 705798
rect 128382 705242 128414 705798
rect 127794 669454 128414 705242
rect 127794 668898 127826 669454
rect 128382 668898 128414 669454
rect 127794 633454 128414 668898
rect 127794 632898 127826 633454
rect 128382 632898 128414 633454
rect 127794 597454 128414 632898
rect 127794 596898 127826 597454
rect 128382 596898 128414 597454
rect 127794 561454 128414 596898
rect 127794 560898 127826 561454
rect 128382 560898 128414 561454
rect 127794 525454 128414 560898
rect 127794 524898 127826 525454
rect 128382 524898 128414 525454
rect 127794 489454 128414 524898
rect 127794 488898 127826 489454
rect 128382 488898 128414 489454
rect 127794 453454 128414 488898
rect 127794 452898 127826 453454
rect 128382 452898 128414 453454
rect 127794 417454 128414 452898
rect 127794 416898 127826 417454
rect 128382 416898 128414 417454
rect 127794 381454 128414 416898
rect 127794 380898 127826 381454
rect 128382 380898 128414 381454
rect 127794 345454 128414 380898
rect 127794 344898 127826 345454
rect 128382 344898 128414 345454
rect 127794 309454 128414 344898
rect 127794 308898 127826 309454
rect 128382 308898 128414 309454
rect 127794 273454 128414 308898
rect 127794 272898 127826 273454
rect 128382 272898 128414 273454
rect 127794 237454 128414 272898
rect 127794 236898 127826 237454
rect 128382 236898 128414 237454
rect 127794 201454 128414 236898
rect 127794 200898 127826 201454
rect 128382 200898 128414 201454
rect 127794 165454 128414 200898
rect 127794 164898 127826 165454
rect 128382 164898 128414 165454
rect 127794 129454 128414 164898
rect 127794 128898 127826 129454
rect 128382 128898 128414 129454
rect 127794 93454 128414 128898
rect 127794 92898 127826 93454
rect 128382 92898 128414 93454
rect 127794 57454 128414 92898
rect 127794 56898 127826 57454
rect 128382 56898 128414 57454
rect 127794 21454 128414 56898
rect 127794 20898 127826 21454
rect 128382 20898 128414 21454
rect 127794 -1306 128414 20898
rect 127794 -1862 127826 -1306
rect 128382 -1862 128414 -1306
rect 127794 -1894 128414 -1862
rect 131514 673174 132134 707162
rect 131514 672618 131546 673174
rect 132102 672618 132134 673174
rect 131514 637174 132134 672618
rect 131514 636618 131546 637174
rect 132102 636618 132134 637174
rect 131514 601174 132134 636618
rect 131514 600618 131546 601174
rect 132102 600618 132134 601174
rect 131514 565174 132134 600618
rect 131514 564618 131546 565174
rect 132102 564618 132134 565174
rect 131514 529174 132134 564618
rect 131514 528618 131546 529174
rect 132102 528618 132134 529174
rect 131514 493174 132134 528618
rect 131514 492618 131546 493174
rect 132102 492618 132134 493174
rect 131514 457174 132134 492618
rect 131514 456618 131546 457174
rect 132102 456618 132134 457174
rect 131514 421174 132134 456618
rect 131514 420618 131546 421174
rect 132102 420618 132134 421174
rect 131514 385174 132134 420618
rect 131514 384618 131546 385174
rect 132102 384618 132134 385174
rect 131514 349174 132134 384618
rect 131514 348618 131546 349174
rect 132102 348618 132134 349174
rect 131514 313174 132134 348618
rect 131514 312618 131546 313174
rect 132102 312618 132134 313174
rect 131514 277174 132134 312618
rect 131514 276618 131546 277174
rect 132102 276618 132134 277174
rect 131514 241174 132134 276618
rect 131514 240618 131546 241174
rect 132102 240618 132134 241174
rect 131514 205174 132134 240618
rect 131514 204618 131546 205174
rect 132102 204618 132134 205174
rect 131514 169174 132134 204618
rect 131514 168618 131546 169174
rect 132102 168618 132134 169174
rect 131514 133174 132134 168618
rect 131514 132618 131546 133174
rect 132102 132618 132134 133174
rect 131514 97174 132134 132618
rect 131514 96618 131546 97174
rect 132102 96618 132134 97174
rect 131514 61174 132134 96618
rect 131514 60618 131546 61174
rect 132102 60618 132134 61174
rect 131514 25174 132134 60618
rect 131514 24618 131546 25174
rect 132102 24618 132134 25174
rect 131514 -3226 132134 24618
rect 131514 -3782 131546 -3226
rect 132102 -3782 132134 -3226
rect 131514 -3814 132134 -3782
rect 135234 676894 135854 709082
rect 135234 676338 135266 676894
rect 135822 676338 135854 676894
rect 135234 640894 135854 676338
rect 135234 640338 135266 640894
rect 135822 640338 135854 640894
rect 135234 604894 135854 640338
rect 135234 604338 135266 604894
rect 135822 604338 135854 604894
rect 135234 568894 135854 604338
rect 135234 568338 135266 568894
rect 135822 568338 135854 568894
rect 135234 532894 135854 568338
rect 135234 532338 135266 532894
rect 135822 532338 135854 532894
rect 135234 496894 135854 532338
rect 135234 496338 135266 496894
rect 135822 496338 135854 496894
rect 135234 460894 135854 496338
rect 135234 460338 135266 460894
rect 135822 460338 135854 460894
rect 135234 424894 135854 460338
rect 135234 424338 135266 424894
rect 135822 424338 135854 424894
rect 135234 388894 135854 424338
rect 135234 388338 135266 388894
rect 135822 388338 135854 388894
rect 135234 352894 135854 388338
rect 135234 352338 135266 352894
rect 135822 352338 135854 352894
rect 135234 316894 135854 352338
rect 135234 316338 135266 316894
rect 135822 316338 135854 316894
rect 135234 280894 135854 316338
rect 135234 280338 135266 280894
rect 135822 280338 135854 280894
rect 135234 244894 135854 280338
rect 135234 244338 135266 244894
rect 135822 244338 135854 244894
rect 135234 208894 135854 244338
rect 135234 208338 135266 208894
rect 135822 208338 135854 208894
rect 135234 172894 135854 208338
rect 135234 172338 135266 172894
rect 135822 172338 135854 172894
rect 135234 136894 135854 172338
rect 135234 136338 135266 136894
rect 135822 136338 135854 136894
rect 135234 100894 135854 136338
rect 135234 100338 135266 100894
rect 135822 100338 135854 100894
rect 135234 64894 135854 100338
rect 135234 64338 135266 64894
rect 135822 64338 135854 64894
rect 135234 28894 135854 64338
rect 135234 28338 135266 28894
rect 135822 28338 135854 28894
rect 135234 -5146 135854 28338
rect 135234 -5702 135266 -5146
rect 135822 -5702 135854 -5146
rect 135234 -5734 135854 -5702
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710042 156986 710598
rect 157542 710042 157574 710598
rect 153234 708678 153854 709670
rect 153234 708122 153266 708678
rect 153822 708122 153854 708678
rect 149514 706758 150134 707750
rect 149514 706202 149546 706758
rect 150102 706202 150134 706758
rect 138954 680058 138986 680614
rect 139542 680058 139574 680614
rect 138954 644614 139574 680058
rect 138954 644058 138986 644614
rect 139542 644058 139574 644614
rect 138954 608614 139574 644058
rect 138954 608058 138986 608614
rect 139542 608058 139574 608614
rect 138954 572614 139574 608058
rect 138954 572058 138986 572614
rect 139542 572058 139574 572614
rect 138954 536614 139574 572058
rect 138954 536058 138986 536614
rect 139542 536058 139574 536614
rect 138954 500614 139574 536058
rect 138954 500058 138986 500614
rect 139542 500058 139574 500614
rect 138954 464614 139574 500058
rect 138954 464058 138986 464614
rect 139542 464058 139574 464614
rect 138954 428614 139574 464058
rect 138954 428058 138986 428614
rect 139542 428058 139574 428614
rect 138954 392614 139574 428058
rect 138954 392058 138986 392614
rect 139542 392058 139574 392614
rect 138954 356614 139574 392058
rect 138954 356058 138986 356614
rect 139542 356058 139574 356614
rect 138954 320614 139574 356058
rect 138954 320058 138986 320614
rect 139542 320058 139574 320614
rect 138954 284614 139574 320058
rect 138954 284058 138986 284614
rect 139542 284058 139574 284614
rect 138954 248614 139574 284058
rect 138954 248058 138986 248614
rect 139542 248058 139574 248614
rect 138954 212614 139574 248058
rect 138954 212058 138986 212614
rect 139542 212058 139574 212614
rect 138954 176614 139574 212058
rect 138954 176058 138986 176614
rect 139542 176058 139574 176614
rect 138954 140614 139574 176058
rect 138954 140058 138986 140614
rect 139542 140058 139574 140614
rect 138954 104614 139574 140058
rect 138954 104058 138986 104614
rect 139542 104058 139574 104614
rect 138954 68614 139574 104058
rect 138954 68058 138986 68614
rect 139542 68058 139574 68614
rect 138954 32614 139574 68058
rect 138954 32058 138986 32614
rect 139542 32058 139574 32614
rect 120954 -6662 120986 -6106
rect 121542 -6662 121574 -6106
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 704838 146414 705830
rect 145794 704282 145826 704838
rect 146382 704282 146414 704838
rect 145794 687454 146414 704282
rect 145794 686898 145826 687454
rect 146382 686898 146414 687454
rect 145794 651454 146414 686898
rect 145794 650898 145826 651454
rect 146382 650898 146414 651454
rect 145794 615454 146414 650898
rect 145794 614898 145826 615454
rect 146382 614898 146414 615454
rect 145794 579454 146414 614898
rect 145794 578898 145826 579454
rect 146382 578898 146414 579454
rect 145794 543454 146414 578898
rect 145794 542898 145826 543454
rect 146382 542898 146414 543454
rect 145794 507454 146414 542898
rect 145794 506898 145826 507454
rect 146382 506898 146414 507454
rect 145794 471454 146414 506898
rect 145794 470898 145826 471454
rect 146382 470898 146414 471454
rect 145794 435454 146414 470898
rect 145794 434898 145826 435454
rect 146382 434898 146414 435454
rect 145794 399454 146414 434898
rect 145794 398898 145826 399454
rect 146382 398898 146414 399454
rect 145794 363454 146414 398898
rect 145794 362898 145826 363454
rect 146382 362898 146414 363454
rect 145794 327454 146414 362898
rect 145794 326898 145826 327454
rect 146382 326898 146414 327454
rect 145794 291454 146414 326898
rect 145794 290898 145826 291454
rect 146382 290898 146414 291454
rect 145794 255454 146414 290898
rect 145794 254898 145826 255454
rect 146382 254898 146414 255454
rect 145794 219454 146414 254898
rect 145794 218898 145826 219454
rect 146382 218898 146414 219454
rect 145794 183454 146414 218898
rect 145794 182898 145826 183454
rect 146382 182898 146414 183454
rect 145794 147454 146414 182898
rect 145794 146898 145826 147454
rect 146382 146898 146414 147454
rect 145794 111454 146414 146898
rect 145794 110898 145826 111454
rect 146382 110898 146414 111454
rect 145794 75454 146414 110898
rect 145794 74898 145826 75454
rect 146382 74898 146414 75454
rect 145794 39454 146414 74898
rect 145794 38898 145826 39454
rect 146382 38898 146414 39454
rect 145794 3454 146414 38898
rect 145794 2898 145826 3454
rect 146382 2898 146414 3454
rect 145794 -346 146414 2898
rect 145794 -902 145826 -346
rect 146382 -902 146414 -346
rect 145794 -1894 146414 -902
rect 149514 691174 150134 706202
rect 149514 690618 149546 691174
rect 150102 690618 150134 691174
rect 149514 655174 150134 690618
rect 149514 654618 149546 655174
rect 150102 654618 150134 655174
rect 149514 619174 150134 654618
rect 149514 618618 149546 619174
rect 150102 618618 150134 619174
rect 149514 583174 150134 618618
rect 149514 582618 149546 583174
rect 150102 582618 150134 583174
rect 149514 547174 150134 582618
rect 149514 546618 149546 547174
rect 150102 546618 150134 547174
rect 149514 511174 150134 546618
rect 149514 510618 149546 511174
rect 150102 510618 150134 511174
rect 149514 475174 150134 510618
rect 149514 474618 149546 475174
rect 150102 474618 150134 475174
rect 149514 439174 150134 474618
rect 149514 438618 149546 439174
rect 150102 438618 150134 439174
rect 149514 403174 150134 438618
rect 149514 402618 149546 403174
rect 150102 402618 150134 403174
rect 149514 367174 150134 402618
rect 149514 366618 149546 367174
rect 150102 366618 150134 367174
rect 149514 331174 150134 366618
rect 149514 330618 149546 331174
rect 150102 330618 150134 331174
rect 149514 295174 150134 330618
rect 149514 294618 149546 295174
rect 150102 294618 150134 295174
rect 149514 259174 150134 294618
rect 149514 258618 149546 259174
rect 150102 258618 150134 259174
rect 149514 223174 150134 258618
rect 149514 222618 149546 223174
rect 150102 222618 150134 223174
rect 149514 187174 150134 222618
rect 149514 186618 149546 187174
rect 150102 186618 150134 187174
rect 149514 151174 150134 186618
rect 149514 150618 149546 151174
rect 150102 150618 150134 151174
rect 149514 115174 150134 150618
rect 149514 114618 149546 115174
rect 150102 114618 150134 115174
rect 149514 79174 150134 114618
rect 149514 78618 149546 79174
rect 150102 78618 150134 79174
rect 149514 43174 150134 78618
rect 149514 42618 149546 43174
rect 150102 42618 150134 43174
rect 149514 7174 150134 42618
rect 149514 6618 149546 7174
rect 150102 6618 150134 7174
rect 149514 -2266 150134 6618
rect 149514 -2822 149546 -2266
rect 150102 -2822 150134 -2266
rect 149514 -3814 150134 -2822
rect 153234 694894 153854 708122
rect 153234 694338 153266 694894
rect 153822 694338 153854 694894
rect 153234 658894 153854 694338
rect 153234 658338 153266 658894
rect 153822 658338 153854 658894
rect 153234 622894 153854 658338
rect 153234 622338 153266 622894
rect 153822 622338 153854 622894
rect 153234 586894 153854 622338
rect 153234 586338 153266 586894
rect 153822 586338 153854 586894
rect 153234 550894 153854 586338
rect 153234 550338 153266 550894
rect 153822 550338 153854 550894
rect 153234 514894 153854 550338
rect 153234 514338 153266 514894
rect 153822 514338 153854 514894
rect 153234 478894 153854 514338
rect 153234 478338 153266 478894
rect 153822 478338 153854 478894
rect 153234 442894 153854 478338
rect 153234 442338 153266 442894
rect 153822 442338 153854 442894
rect 153234 406894 153854 442338
rect 153234 406338 153266 406894
rect 153822 406338 153854 406894
rect 153234 370894 153854 406338
rect 153234 370338 153266 370894
rect 153822 370338 153854 370894
rect 153234 334894 153854 370338
rect 153234 334338 153266 334894
rect 153822 334338 153854 334894
rect 153234 298894 153854 334338
rect 153234 298338 153266 298894
rect 153822 298338 153854 298894
rect 153234 262894 153854 298338
rect 153234 262338 153266 262894
rect 153822 262338 153854 262894
rect 153234 226894 153854 262338
rect 153234 226338 153266 226894
rect 153822 226338 153854 226894
rect 153234 190894 153854 226338
rect 153234 190338 153266 190894
rect 153822 190338 153854 190894
rect 153234 154894 153854 190338
rect 153234 154338 153266 154894
rect 153822 154338 153854 154894
rect 153234 118894 153854 154338
rect 153234 118338 153266 118894
rect 153822 118338 153854 118894
rect 153234 82894 153854 118338
rect 153234 82338 153266 82894
rect 153822 82338 153854 82894
rect 153234 46894 153854 82338
rect 153234 46338 153266 46894
rect 153822 46338 153854 46894
rect 153234 10894 153854 46338
rect 153234 10338 153266 10894
rect 153822 10338 153854 10894
rect 153234 -4186 153854 10338
rect 153234 -4742 153266 -4186
rect 153822 -4742 153854 -4186
rect 153234 -5734 153854 -4742
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711002 174986 711558
rect 175542 711002 175574 711558
rect 171234 709638 171854 709670
rect 171234 709082 171266 709638
rect 171822 709082 171854 709638
rect 167514 707718 168134 707750
rect 167514 707162 167546 707718
rect 168102 707162 168134 707718
rect 156954 698058 156986 698614
rect 157542 698058 157574 698614
rect 156954 662614 157574 698058
rect 156954 662058 156986 662614
rect 157542 662058 157574 662614
rect 156954 626614 157574 662058
rect 156954 626058 156986 626614
rect 157542 626058 157574 626614
rect 156954 590614 157574 626058
rect 156954 590058 156986 590614
rect 157542 590058 157574 590614
rect 156954 554614 157574 590058
rect 156954 554058 156986 554614
rect 157542 554058 157574 554614
rect 156954 518614 157574 554058
rect 156954 518058 156986 518614
rect 157542 518058 157574 518614
rect 156954 482614 157574 518058
rect 156954 482058 156986 482614
rect 157542 482058 157574 482614
rect 156954 446614 157574 482058
rect 156954 446058 156986 446614
rect 157542 446058 157574 446614
rect 156954 410614 157574 446058
rect 156954 410058 156986 410614
rect 157542 410058 157574 410614
rect 156954 374614 157574 410058
rect 156954 374058 156986 374614
rect 157542 374058 157574 374614
rect 156954 338614 157574 374058
rect 156954 338058 156986 338614
rect 157542 338058 157574 338614
rect 156954 302614 157574 338058
rect 156954 302058 156986 302614
rect 157542 302058 157574 302614
rect 156954 266614 157574 302058
rect 156954 266058 156986 266614
rect 157542 266058 157574 266614
rect 156954 230614 157574 266058
rect 156954 230058 156986 230614
rect 157542 230058 157574 230614
rect 156954 194614 157574 230058
rect 156954 194058 156986 194614
rect 157542 194058 157574 194614
rect 156954 158614 157574 194058
rect 156954 158058 156986 158614
rect 157542 158058 157574 158614
rect 156954 122614 157574 158058
rect 156954 122058 156986 122614
rect 157542 122058 157574 122614
rect 156954 86614 157574 122058
rect 156954 86058 156986 86614
rect 157542 86058 157574 86614
rect 156954 50614 157574 86058
rect 156954 50058 156986 50614
rect 157542 50058 157574 50614
rect 156954 14614 157574 50058
rect 156954 14058 156986 14614
rect 157542 14058 157574 14614
rect 138954 -7622 138986 -7066
rect 139542 -7622 139574 -7066
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 705798 164414 705830
rect 163794 705242 163826 705798
rect 164382 705242 164414 705798
rect 163794 669454 164414 705242
rect 163794 668898 163826 669454
rect 164382 668898 164414 669454
rect 163794 633454 164414 668898
rect 163794 632898 163826 633454
rect 164382 632898 164414 633454
rect 163794 597454 164414 632898
rect 163794 596898 163826 597454
rect 164382 596898 164414 597454
rect 163794 561454 164414 596898
rect 163794 560898 163826 561454
rect 164382 560898 164414 561454
rect 163794 525454 164414 560898
rect 163794 524898 163826 525454
rect 164382 524898 164414 525454
rect 163794 489454 164414 524898
rect 163794 488898 163826 489454
rect 164382 488898 164414 489454
rect 163794 453454 164414 488898
rect 163794 452898 163826 453454
rect 164382 452898 164414 453454
rect 163794 417454 164414 452898
rect 163794 416898 163826 417454
rect 164382 416898 164414 417454
rect 163794 381454 164414 416898
rect 163794 380898 163826 381454
rect 164382 380898 164414 381454
rect 163794 345454 164414 380898
rect 163794 344898 163826 345454
rect 164382 344898 164414 345454
rect 163794 309454 164414 344898
rect 163794 308898 163826 309454
rect 164382 308898 164414 309454
rect 163794 273454 164414 308898
rect 163794 272898 163826 273454
rect 164382 272898 164414 273454
rect 163794 237454 164414 272898
rect 163794 236898 163826 237454
rect 164382 236898 164414 237454
rect 163794 201454 164414 236898
rect 163794 200898 163826 201454
rect 164382 200898 164414 201454
rect 163794 165454 164414 200898
rect 163794 164898 163826 165454
rect 164382 164898 164414 165454
rect 163794 129454 164414 164898
rect 163794 128898 163826 129454
rect 164382 128898 164414 129454
rect 163794 93454 164414 128898
rect 163794 92898 163826 93454
rect 164382 92898 164414 93454
rect 163794 57454 164414 92898
rect 163794 56898 163826 57454
rect 164382 56898 164414 57454
rect 163794 21454 164414 56898
rect 163794 20898 163826 21454
rect 164382 20898 164414 21454
rect 163794 -1306 164414 20898
rect 163794 -1862 163826 -1306
rect 164382 -1862 164414 -1306
rect 163794 -1894 164414 -1862
rect 167514 673174 168134 707162
rect 167514 672618 167546 673174
rect 168102 672618 168134 673174
rect 167514 637174 168134 672618
rect 167514 636618 167546 637174
rect 168102 636618 168134 637174
rect 167514 601174 168134 636618
rect 167514 600618 167546 601174
rect 168102 600618 168134 601174
rect 167514 565174 168134 600618
rect 167514 564618 167546 565174
rect 168102 564618 168134 565174
rect 167514 529174 168134 564618
rect 167514 528618 167546 529174
rect 168102 528618 168134 529174
rect 167514 493174 168134 528618
rect 167514 492618 167546 493174
rect 168102 492618 168134 493174
rect 167514 457174 168134 492618
rect 167514 456618 167546 457174
rect 168102 456618 168134 457174
rect 167514 421174 168134 456618
rect 167514 420618 167546 421174
rect 168102 420618 168134 421174
rect 167514 385174 168134 420618
rect 167514 384618 167546 385174
rect 168102 384618 168134 385174
rect 167514 349174 168134 384618
rect 167514 348618 167546 349174
rect 168102 348618 168134 349174
rect 167514 313174 168134 348618
rect 167514 312618 167546 313174
rect 168102 312618 168134 313174
rect 167514 277174 168134 312618
rect 167514 276618 167546 277174
rect 168102 276618 168134 277174
rect 167514 241174 168134 276618
rect 167514 240618 167546 241174
rect 168102 240618 168134 241174
rect 167514 205174 168134 240618
rect 167514 204618 167546 205174
rect 168102 204618 168134 205174
rect 167514 169174 168134 204618
rect 167514 168618 167546 169174
rect 168102 168618 168134 169174
rect 167514 133174 168134 168618
rect 167514 132618 167546 133174
rect 168102 132618 168134 133174
rect 167514 97174 168134 132618
rect 167514 96618 167546 97174
rect 168102 96618 168134 97174
rect 167514 61174 168134 96618
rect 167514 60618 167546 61174
rect 168102 60618 168134 61174
rect 167514 25174 168134 60618
rect 167514 24618 167546 25174
rect 168102 24618 168134 25174
rect 167514 -3226 168134 24618
rect 167514 -3782 167546 -3226
rect 168102 -3782 168134 -3226
rect 167514 -3814 168134 -3782
rect 171234 676894 171854 709082
rect 171234 676338 171266 676894
rect 171822 676338 171854 676894
rect 171234 640894 171854 676338
rect 171234 640338 171266 640894
rect 171822 640338 171854 640894
rect 171234 604894 171854 640338
rect 171234 604338 171266 604894
rect 171822 604338 171854 604894
rect 171234 568894 171854 604338
rect 171234 568338 171266 568894
rect 171822 568338 171854 568894
rect 171234 532894 171854 568338
rect 171234 532338 171266 532894
rect 171822 532338 171854 532894
rect 171234 496894 171854 532338
rect 171234 496338 171266 496894
rect 171822 496338 171854 496894
rect 171234 460894 171854 496338
rect 171234 460338 171266 460894
rect 171822 460338 171854 460894
rect 171234 424894 171854 460338
rect 171234 424338 171266 424894
rect 171822 424338 171854 424894
rect 171234 388894 171854 424338
rect 171234 388338 171266 388894
rect 171822 388338 171854 388894
rect 171234 352894 171854 388338
rect 171234 352338 171266 352894
rect 171822 352338 171854 352894
rect 171234 316894 171854 352338
rect 171234 316338 171266 316894
rect 171822 316338 171854 316894
rect 171234 280894 171854 316338
rect 171234 280338 171266 280894
rect 171822 280338 171854 280894
rect 171234 244894 171854 280338
rect 171234 244338 171266 244894
rect 171822 244338 171854 244894
rect 171234 208894 171854 244338
rect 171234 208338 171266 208894
rect 171822 208338 171854 208894
rect 171234 172894 171854 208338
rect 171234 172338 171266 172894
rect 171822 172338 171854 172894
rect 171234 136894 171854 172338
rect 171234 136338 171266 136894
rect 171822 136338 171854 136894
rect 171234 100894 171854 136338
rect 171234 100338 171266 100894
rect 171822 100338 171854 100894
rect 171234 64894 171854 100338
rect 171234 64338 171266 64894
rect 171822 64338 171854 64894
rect 171234 28894 171854 64338
rect 171234 28338 171266 28894
rect 171822 28338 171854 28894
rect 171234 -5146 171854 28338
rect 171234 -5702 171266 -5146
rect 171822 -5702 171854 -5146
rect 171234 -5734 171854 -5702
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710042 192986 710598
rect 193542 710042 193574 710598
rect 189234 708678 189854 709670
rect 189234 708122 189266 708678
rect 189822 708122 189854 708678
rect 185514 706758 186134 707750
rect 185514 706202 185546 706758
rect 186102 706202 186134 706758
rect 174954 680058 174986 680614
rect 175542 680058 175574 680614
rect 174954 644614 175574 680058
rect 174954 644058 174986 644614
rect 175542 644058 175574 644614
rect 174954 608614 175574 644058
rect 174954 608058 174986 608614
rect 175542 608058 175574 608614
rect 174954 572614 175574 608058
rect 174954 572058 174986 572614
rect 175542 572058 175574 572614
rect 174954 536614 175574 572058
rect 174954 536058 174986 536614
rect 175542 536058 175574 536614
rect 174954 500614 175574 536058
rect 174954 500058 174986 500614
rect 175542 500058 175574 500614
rect 174954 464614 175574 500058
rect 174954 464058 174986 464614
rect 175542 464058 175574 464614
rect 174954 428614 175574 464058
rect 174954 428058 174986 428614
rect 175542 428058 175574 428614
rect 174954 392614 175574 428058
rect 174954 392058 174986 392614
rect 175542 392058 175574 392614
rect 174954 356614 175574 392058
rect 174954 356058 174986 356614
rect 175542 356058 175574 356614
rect 174954 320614 175574 356058
rect 174954 320058 174986 320614
rect 175542 320058 175574 320614
rect 174954 284614 175574 320058
rect 174954 284058 174986 284614
rect 175542 284058 175574 284614
rect 174954 248614 175574 284058
rect 174954 248058 174986 248614
rect 175542 248058 175574 248614
rect 174954 212614 175574 248058
rect 174954 212058 174986 212614
rect 175542 212058 175574 212614
rect 174954 176614 175574 212058
rect 174954 176058 174986 176614
rect 175542 176058 175574 176614
rect 174954 140614 175574 176058
rect 174954 140058 174986 140614
rect 175542 140058 175574 140614
rect 174954 104614 175574 140058
rect 174954 104058 174986 104614
rect 175542 104058 175574 104614
rect 174954 68614 175574 104058
rect 174954 68058 174986 68614
rect 175542 68058 175574 68614
rect 174954 32614 175574 68058
rect 174954 32058 174986 32614
rect 175542 32058 175574 32614
rect 156954 -6662 156986 -6106
rect 157542 -6662 157574 -6106
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 704838 182414 705830
rect 181794 704282 181826 704838
rect 182382 704282 182414 704838
rect 181794 687454 182414 704282
rect 181794 686898 181826 687454
rect 182382 686898 182414 687454
rect 181794 651454 182414 686898
rect 181794 650898 181826 651454
rect 182382 650898 182414 651454
rect 181794 615454 182414 650898
rect 181794 614898 181826 615454
rect 182382 614898 182414 615454
rect 181794 579454 182414 614898
rect 181794 578898 181826 579454
rect 182382 578898 182414 579454
rect 181794 543454 182414 578898
rect 181794 542898 181826 543454
rect 182382 542898 182414 543454
rect 181794 507454 182414 542898
rect 181794 506898 181826 507454
rect 182382 506898 182414 507454
rect 181794 471454 182414 506898
rect 181794 470898 181826 471454
rect 182382 470898 182414 471454
rect 181794 435454 182414 470898
rect 181794 434898 181826 435454
rect 182382 434898 182414 435454
rect 181794 399454 182414 434898
rect 181794 398898 181826 399454
rect 182382 398898 182414 399454
rect 181794 363454 182414 398898
rect 181794 362898 181826 363454
rect 182382 362898 182414 363454
rect 181794 327454 182414 362898
rect 181794 326898 181826 327454
rect 182382 326898 182414 327454
rect 181794 291454 182414 326898
rect 181794 290898 181826 291454
rect 182382 290898 182414 291454
rect 181794 255454 182414 290898
rect 181794 254898 181826 255454
rect 182382 254898 182414 255454
rect 181794 219454 182414 254898
rect 181794 218898 181826 219454
rect 182382 218898 182414 219454
rect 181794 183454 182414 218898
rect 181794 182898 181826 183454
rect 182382 182898 182414 183454
rect 181794 147454 182414 182898
rect 181794 146898 181826 147454
rect 182382 146898 182414 147454
rect 181794 111454 182414 146898
rect 181794 110898 181826 111454
rect 182382 110898 182414 111454
rect 181794 75454 182414 110898
rect 181794 74898 181826 75454
rect 182382 74898 182414 75454
rect 181794 39454 182414 74898
rect 181794 38898 181826 39454
rect 182382 38898 182414 39454
rect 181794 3454 182414 38898
rect 181794 2898 181826 3454
rect 182382 2898 182414 3454
rect 181794 -346 182414 2898
rect 181794 -902 181826 -346
rect 182382 -902 182414 -346
rect 181794 -1894 182414 -902
rect 185514 691174 186134 706202
rect 185514 690618 185546 691174
rect 186102 690618 186134 691174
rect 185514 655174 186134 690618
rect 185514 654618 185546 655174
rect 186102 654618 186134 655174
rect 185514 619174 186134 654618
rect 185514 618618 185546 619174
rect 186102 618618 186134 619174
rect 185514 583174 186134 618618
rect 185514 582618 185546 583174
rect 186102 582618 186134 583174
rect 185514 547174 186134 582618
rect 185514 546618 185546 547174
rect 186102 546618 186134 547174
rect 185514 511174 186134 546618
rect 185514 510618 185546 511174
rect 186102 510618 186134 511174
rect 185514 475174 186134 510618
rect 185514 474618 185546 475174
rect 186102 474618 186134 475174
rect 185514 439174 186134 474618
rect 185514 438618 185546 439174
rect 186102 438618 186134 439174
rect 185514 403174 186134 438618
rect 185514 402618 185546 403174
rect 186102 402618 186134 403174
rect 185514 367174 186134 402618
rect 185514 366618 185546 367174
rect 186102 366618 186134 367174
rect 185514 331174 186134 366618
rect 185514 330618 185546 331174
rect 186102 330618 186134 331174
rect 185514 295174 186134 330618
rect 185514 294618 185546 295174
rect 186102 294618 186134 295174
rect 185514 259174 186134 294618
rect 185514 258618 185546 259174
rect 186102 258618 186134 259174
rect 185514 223174 186134 258618
rect 185514 222618 185546 223174
rect 186102 222618 186134 223174
rect 185514 187174 186134 222618
rect 185514 186618 185546 187174
rect 186102 186618 186134 187174
rect 185514 151174 186134 186618
rect 185514 150618 185546 151174
rect 186102 150618 186134 151174
rect 185514 115174 186134 150618
rect 185514 114618 185546 115174
rect 186102 114618 186134 115174
rect 185514 79174 186134 114618
rect 185514 78618 185546 79174
rect 186102 78618 186134 79174
rect 185514 43174 186134 78618
rect 185514 42618 185546 43174
rect 186102 42618 186134 43174
rect 185514 7174 186134 42618
rect 185514 6618 185546 7174
rect 186102 6618 186134 7174
rect 185514 -2266 186134 6618
rect 185514 -2822 185546 -2266
rect 186102 -2822 186134 -2266
rect 185514 -3814 186134 -2822
rect 189234 694894 189854 708122
rect 189234 694338 189266 694894
rect 189822 694338 189854 694894
rect 189234 658894 189854 694338
rect 189234 658338 189266 658894
rect 189822 658338 189854 658894
rect 189234 622894 189854 658338
rect 189234 622338 189266 622894
rect 189822 622338 189854 622894
rect 189234 586894 189854 622338
rect 189234 586338 189266 586894
rect 189822 586338 189854 586894
rect 189234 550894 189854 586338
rect 189234 550338 189266 550894
rect 189822 550338 189854 550894
rect 189234 514894 189854 550338
rect 189234 514338 189266 514894
rect 189822 514338 189854 514894
rect 189234 478894 189854 514338
rect 189234 478338 189266 478894
rect 189822 478338 189854 478894
rect 189234 442894 189854 478338
rect 189234 442338 189266 442894
rect 189822 442338 189854 442894
rect 189234 406894 189854 442338
rect 189234 406338 189266 406894
rect 189822 406338 189854 406894
rect 189234 370894 189854 406338
rect 189234 370338 189266 370894
rect 189822 370338 189854 370894
rect 189234 334894 189854 370338
rect 189234 334338 189266 334894
rect 189822 334338 189854 334894
rect 189234 298894 189854 334338
rect 189234 298338 189266 298894
rect 189822 298338 189854 298894
rect 189234 262894 189854 298338
rect 189234 262338 189266 262894
rect 189822 262338 189854 262894
rect 189234 226894 189854 262338
rect 189234 226338 189266 226894
rect 189822 226338 189854 226894
rect 189234 190894 189854 226338
rect 189234 190338 189266 190894
rect 189822 190338 189854 190894
rect 189234 154894 189854 190338
rect 189234 154338 189266 154894
rect 189822 154338 189854 154894
rect 189234 118894 189854 154338
rect 189234 118338 189266 118894
rect 189822 118338 189854 118894
rect 189234 82894 189854 118338
rect 189234 82338 189266 82894
rect 189822 82338 189854 82894
rect 189234 46894 189854 82338
rect 189234 46338 189266 46894
rect 189822 46338 189854 46894
rect 189234 10894 189854 46338
rect 189234 10338 189266 10894
rect 189822 10338 189854 10894
rect 189234 -4186 189854 10338
rect 189234 -4742 189266 -4186
rect 189822 -4742 189854 -4186
rect 189234 -5734 189854 -4742
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711002 210986 711558
rect 211542 711002 211574 711558
rect 207234 709638 207854 709670
rect 207234 709082 207266 709638
rect 207822 709082 207854 709638
rect 203514 707718 204134 707750
rect 203514 707162 203546 707718
rect 204102 707162 204134 707718
rect 192954 698058 192986 698614
rect 193542 698058 193574 698614
rect 192954 662614 193574 698058
rect 192954 662058 192986 662614
rect 193542 662058 193574 662614
rect 192954 626614 193574 662058
rect 192954 626058 192986 626614
rect 193542 626058 193574 626614
rect 192954 590614 193574 626058
rect 192954 590058 192986 590614
rect 193542 590058 193574 590614
rect 192954 554614 193574 590058
rect 192954 554058 192986 554614
rect 193542 554058 193574 554614
rect 192954 518614 193574 554058
rect 192954 518058 192986 518614
rect 193542 518058 193574 518614
rect 192954 482614 193574 518058
rect 192954 482058 192986 482614
rect 193542 482058 193574 482614
rect 192954 446614 193574 482058
rect 192954 446058 192986 446614
rect 193542 446058 193574 446614
rect 192954 410614 193574 446058
rect 192954 410058 192986 410614
rect 193542 410058 193574 410614
rect 192954 374614 193574 410058
rect 192954 374058 192986 374614
rect 193542 374058 193574 374614
rect 192954 338614 193574 374058
rect 192954 338058 192986 338614
rect 193542 338058 193574 338614
rect 192954 302614 193574 338058
rect 192954 302058 192986 302614
rect 193542 302058 193574 302614
rect 192954 266614 193574 302058
rect 192954 266058 192986 266614
rect 193542 266058 193574 266614
rect 192954 230614 193574 266058
rect 192954 230058 192986 230614
rect 193542 230058 193574 230614
rect 192954 194614 193574 230058
rect 192954 194058 192986 194614
rect 193542 194058 193574 194614
rect 192954 158614 193574 194058
rect 192954 158058 192986 158614
rect 193542 158058 193574 158614
rect 192954 122614 193574 158058
rect 192954 122058 192986 122614
rect 193542 122058 193574 122614
rect 192954 86614 193574 122058
rect 192954 86058 192986 86614
rect 193542 86058 193574 86614
rect 192954 50614 193574 86058
rect 192954 50058 192986 50614
rect 193542 50058 193574 50614
rect 192954 14614 193574 50058
rect 192954 14058 192986 14614
rect 193542 14058 193574 14614
rect 174954 -7622 174986 -7066
rect 175542 -7622 175574 -7066
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 705798 200414 705830
rect 199794 705242 199826 705798
rect 200382 705242 200414 705798
rect 199794 669454 200414 705242
rect 199794 668898 199826 669454
rect 200382 668898 200414 669454
rect 199794 633454 200414 668898
rect 199794 632898 199826 633454
rect 200382 632898 200414 633454
rect 199794 597454 200414 632898
rect 199794 596898 199826 597454
rect 200382 596898 200414 597454
rect 199794 561454 200414 596898
rect 199794 560898 199826 561454
rect 200382 560898 200414 561454
rect 199794 525454 200414 560898
rect 199794 524898 199826 525454
rect 200382 524898 200414 525454
rect 199794 489454 200414 524898
rect 199794 488898 199826 489454
rect 200382 488898 200414 489454
rect 199794 453454 200414 488898
rect 199794 452898 199826 453454
rect 200382 452898 200414 453454
rect 199794 417454 200414 452898
rect 199794 416898 199826 417454
rect 200382 416898 200414 417454
rect 199794 381454 200414 416898
rect 199794 380898 199826 381454
rect 200382 380898 200414 381454
rect 199794 345454 200414 380898
rect 199794 344898 199826 345454
rect 200382 344898 200414 345454
rect 199794 309454 200414 344898
rect 199794 308898 199826 309454
rect 200382 308898 200414 309454
rect 199794 273454 200414 308898
rect 199794 272898 199826 273454
rect 200382 272898 200414 273454
rect 199794 237454 200414 272898
rect 199794 236898 199826 237454
rect 200382 236898 200414 237454
rect 199794 201454 200414 236898
rect 199794 200898 199826 201454
rect 200382 200898 200414 201454
rect 199794 165454 200414 200898
rect 199794 164898 199826 165454
rect 200382 164898 200414 165454
rect 199794 129454 200414 164898
rect 199794 128898 199826 129454
rect 200382 128898 200414 129454
rect 199794 93454 200414 128898
rect 199794 92898 199826 93454
rect 200382 92898 200414 93454
rect 199794 57454 200414 92898
rect 199794 56898 199826 57454
rect 200382 56898 200414 57454
rect 199794 21454 200414 56898
rect 199794 20898 199826 21454
rect 200382 20898 200414 21454
rect 199794 -1306 200414 20898
rect 199794 -1862 199826 -1306
rect 200382 -1862 200414 -1306
rect 199794 -1894 200414 -1862
rect 203514 673174 204134 707162
rect 203514 672618 203546 673174
rect 204102 672618 204134 673174
rect 203514 637174 204134 672618
rect 203514 636618 203546 637174
rect 204102 636618 204134 637174
rect 203514 601174 204134 636618
rect 203514 600618 203546 601174
rect 204102 600618 204134 601174
rect 203514 565174 204134 600618
rect 203514 564618 203546 565174
rect 204102 564618 204134 565174
rect 203514 529174 204134 564618
rect 203514 528618 203546 529174
rect 204102 528618 204134 529174
rect 203514 493174 204134 528618
rect 203514 492618 203546 493174
rect 204102 492618 204134 493174
rect 203514 457174 204134 492618
rect 203514 456618 203546 457174
rect 204102 456618 204134 457174
rect 203514 421174 204134 456618
rect 203514 420618 203546 421174
rect 204102 420618 204134 421174
rect 203514 385174 204134 420618
rect 203514 384618 203546 385174
rect 204102 384618 204134 385174
rect 203514 349174 204134 384618
rect 203514 348618 203546 349174
rect 204102 348618 204134 349174
rect 203514 313174 204134 348618
rect 203514 312618 203546 313174
rect 204102 312618 204134 313174
rect 203514 277174 204134 312618
rect 203514 276618 203546 277174
rect 204102 276618 204134 277174
rect 203514 241174 204134 276618
rect 203514 240618 203546 241174
rect 204102 240618 204134 241174
rect 203514 205174 204134 240618
rect 203514 204618 203546 205174
rect 204102 204618 204134 205174
rect 203514 169174 204134 204618
rect 203514 168618 203546 169174
rect 204102 168618 204134 169174
rect 203514 133174 204134 168618
rect 203514 132618 203546 133174
rect 204102 132618 204134 133174
rect 203514 97174 204134 132618
rect 203514 96618 203546 97174
rect 204102 96618 204134 97174
rect 203514 61174 204134 96618
rect 203514 60618 203546 61174
rect 204102 60618 204134 61174
rect 203514 25174 204134 60618
rect 203514 24618 203546 25174
rect 204102 24618 204134 25174
rect 203514 -3226 204134 24618
rect 203514 -3782 203546 -3226
rect 204102 -3782 204134 -3226
rect 203514 -3814 204134 -3782
rect 207234 676894 207854 709082
rect 207234 676338 207266 676894
rect 207822 676338 207854 676894
rect 207234 640894 207854 676338
rect 207234 640338 207266 640894
rect 207822 640338 207854 640894
rect 207234 604894 207854 640338
rect 207234 604338 207266 604894
rect 207822 604338 207854 604894
rect 207234 568894 207854 604338
rect 207234 568338 207266 568894
rect 207822 568338 207854 568894
rect 207234 532894 207854 568338
rect 207234 532338 207266 532894
rect 207822 532338 207854 532894
rect 207234 496894 207854 532338
rect 207234 496338 207266 496894
rect 207822 496338 207854 496894
rect 207234 460894 207854 496338
rect 207234 460338 207266 460894
rect 207822 460338 207854 460894
rect 207234 424894 207854 460338
rect 207234 424338 207266 424894
rect 207822 424338 207854 424894
rect 207234 388894 207854 424338
rect 207234 388338 207266 388894
rect 207822 388338 207854 388894
rect 207234 352894 207854 388338
rect 207234 352338 207266 352894
rect 207822 352338 207854 352894
rect 207234 316894 207854 352338
rect 207234 316338 207266 316894
rect 207822 316338 207854 316894
rect 207234 280894 207854 316338
rect 207234 280338 207266 280894
rect 207822 280338 207854 280894
rect 207234 244894 207854 280338
rect 207234 244338 207266 244894
rect 207822 244338 207854 244894
rect 207234 208894 207854 244338
rect 207234 208338 207266 208894
rect 207822 208338 207854 208894
rect 207234 172894 207854 208338
rect 207234 172338 207266 172894
rect 207822 172338 207854 172894
rect 207234 136894 207854 172338
rect 207234 136338 207266 136894
rect 207822 136338 207854 136894
rect 207234 100894 207854 136338
rect 207234 100338 207266 100894
rect 207822 100338 207854 100894
rect 207234 64894 207854 100338
rect 207234 64338 207266 64894
rect 207822 64338 207854 64894
rect 207234 28894 207854 64338
rect 207234 28338 207266 28894
rect 207822 28338 207854 28894
rect 207234 -5146 207854 28338
rect 207234 -5702 207266 -5146
rect 207822 -5702 207854 -5146
rect 207234 -5734 207854 -5702
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710042 228986 710598
rect 229542 710042 229574 710598
rect 225234 708678 225854 709670
rect 225234 708122 225266 708678
rect 225822 708122 225854 708678
rect 221514 706758 222134 707750
rect 221514 706202 221546 706758
rect 222102 706202 222134 706758
rect 210954 680058 210986 680614
rect 211542 680058 211574 680614
rect 210954 644614 211574 680058
rect 210954 644058 210986 644614
rect 211542 644058 211574 644614
rect 210954 608614 211574 644058
rect 210954 608058 210986 608614
rect 211542 608058 211574 608614
rect 210954 572614 211574 608058
rect 210954 572058 210986 572614
rect 211542 572058 211574 572614
rect 210954 536614 211574 572058
rect 210954 536058 210986 536614
rect 211542 536058 211574 536614
rect 210954 500614 211574 536058
rect 210954 500058 210986 500614
rect 211542 500058 211574 500614
rect 210954 464614 211574 500058
rect 210954 464058 210986 464614
rect 211542 464058 211574 464614
rect 210954 428614 211574 464058
rect 210954 428058 210986 428614
rect 211542 428058 211574 428614
rect 210954 392614 211574 428058
rect 210954 392058 210986 392614
rect 211542 392058 211574 392614
rect 210954 356614 211574 392058
rect 210954 356058 210986 356614
rect 211542 356058 211574 356614
rect 210954 320614 211574 356058
rect 210954 320058 210986 320614
rect 211542 320058 211574 320614
rect 210954 284614 211574 320058
rect 210954 284058 210986 284614
rect 211542 284058 211574 284614
rect 210954 248614 211574 284058
rect 210954 248058 210986 248614
rect 211542 248058 211574 248614
rect 210954 212614 211574 248058
rect 210954 212058 210986 212614
rect 211542 212058 211574 212614
rect 210954 176614 211574 212058
rect 210954 176058 210986 176614
rect 211542 176058 211574 176614
rect 210954 140614 211574 176058
rect 210954 140058 210986 140614
rect 211542 140058 211574 140614
rect 210954 104614 211574 140058
rect 210954 104058 210986 104614
rect 211542 104058 211574 104614
rect 210954 68614 211574 104058
rect 210954 68058 210986 68614
rect 211542 68058 211574 68614
rect 210954 32614 211574 68058
rect 210954 32058 210986 32614
rect 211542 32058 211574 32614
rect 192954 -6662 192986 -6106
rect 193542 -6662 193574 -6106
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 704838 218414 705830
rect 217794 704282 217826 704838
rect 218382 704282 218414 704838
rect 217794 687454 218414 704282
rect 217794 686898 217826 687454
rect 218382 686898 218414 687454
rect 217794 651454 218414 686898
rect 217794 650898 217826 651454
rect 218382 650898 218414 651454
rect 217794 615454 218414 650898
rect 217794 614898 217826 615454
rect 218382 614898 218414 615454
rect 217794 579454 218414 614898
rect 217794 578898 217826 579454
rect 218382 578898 218414 579454
rect 217794 543454 218414 578898
rect 217794 542898 217826 543454
rect 218382 542898 218414 543454
rect 217794 507454 218414 542898
rect 217794 506898 217826 507454
rect 218382 506898 218414 507454
rect 217794 471454 218414 506898
rect 217794 470898 217826 471454
rect 218382 470898 218414 471454
rect 217794 435454 218414 470898
rect 217794 434898 217826 435454
rect 218382 434898 218414 435454
rect 217794 399454 218414 434898
rect 217794 398898 217826 399454
rect 218382 398898 218414 399454
rect 217794 363454 218414 398898
rect 217794 362898 217826 363454
rect 218382 362898 218414 363454
rect 217794 327454 218414 362898
rect 217794 326898 217826 327454
rect 218382 326898 218414 327454
rect 217794 291454 218414 326898
rect 217794 290898 217826 291454
rect 218382 290898 218414 291454
rect 217794 255454 218414 290898
rect 217794 254898 217826 255454
rect 218382 254898 218414 255454
rect 217794 219454 218414 254898
rect 217794 218898 217826 219454
rect 218382 218898 218414 219454
rect 217794 183454 218414 218898
rect 217794 182898 217826 183454
rect 218382 182898 218414 183454
rect 217794 147454 218414 182898
rect 217794 146898 217826 147454
rect 218382 146898 218414 147454
rect 217794 111454 218414 146898
rect 217794 110898 217826 111454
rect 218382 110898 218414 111454
rect 217794 75454 218414 110898
rect 217794 74898 217826 75454
rect 218382 74898 218414 75454
rect 217794 39454 218414 74898
rect 217794 38898 217826 39454
rect 218382 38898 218414 39454
rect 217794 3454 218414 38898
rect 217794 2898 217826 3454
rect 218382 2898 218414 3454
rect 217794 -346 218414 2898
rect 217794 -902 217826 -346
rect 218382 -902 218414 -346
rect 217794 -1894 218414 -902
rect 221514 691174 222134 706202
rect 221514 690618 221546 691174
rect 222102 690618 222134 691174
rect 221514 655174 222134 690618
rect 221514 654618 221546 655174
rect 222102 654618 222134 655174
rect 221514 619174 222134 654618
rect 221514 618618 221546 619174
rect 222102 618618 222134 619174
rect 221514 583174 222134 618618
rect 221514 582618 221546 583174
rect 222102 582618 222134 583174
rect 221514 547174 222134 582618
rect 221514 546618 221546 547174
rect 222102 546618 222134 547174
rect 221514 511174 222134 546618
rect 221514 510618 221546 511174
rect 222102 510618 222134 511174
rect 221514 475174 222134 510618
rect 221514 474618 221546 475174
rect 222102 474618 222134 475174
rect 221514 439174 222134 474618
rect 221514 438618 221546 439174
rect 222102 438618 222134 439174
rect 221514 403174 222134 438618
rect 221514 402618 221546 403174
rect 222102 402618 222134 403174
rect 221514 367174 222134 402618
rect 221514 366618 221546 367174
rect 222102 366618 222134 367174
rect 221514 331174 222134 366618
rect 221514 330618 221546 331174
rect 222102 330618 222134 331174
rect 221514 295174 222134 330618
rect 221514 294618 221546 295174
rect 222102 294618 222134 295174
rect 221514 259174 222134 294618
rect 221514 258618 221546 259174
rect 222102 258618 222134 259174
rect 221514 223174 222134 258618
rect 221514 222618 221546 223174
rect 222102 222618 222134 223174
rect 221514 187174 222134 222618
rect 221514 186618 221546 187174
rect 222102 186618 222134 187174
rect 221514 151174 222134 186618
rect 221514 150618 221546 151174
rect 222102 150618 222134 151174
rect 221514 115174 222134 150618
rect 221514 114618 221546 115174
rect 222102 114618 222134 115174
rect 221514 79174 222134 114618
rect 221514 78618 221546 79174
rect 222102 78618 222134 79174
rect 221514 43174 222134 78618
rect 221514 42618 221546 43174
rect 222102 42618 222134 43174
rect 221514 7174 222134 42618
rect 221514 6618 221546 7174
rect 222102 6618 222134 7174
rect 221514 -2266 222134 6618
rect 221514 -2822 221546 -2266
rect 222102 -2822 222134 -2266
rect 221514 -3814 222134 -2822
rect 225234 694894 225854 708122
rect 225234 694338 225266 694894
rect 225822 694338 225854 694894
rect 225234 658894 225854 694338
rect 225234 658338 225266 658894
rect 225822 658338 225854 658894
rect 225234 622894 225854 658338
rect 225234 622338 225266 622894
rect 225822 622338 225854 622894
rect 225234 586894 225854 622338
rect 225234 586338 225266 586894
rect 225822 586338 225854 586894
rect 225234 550894 225854 586338
rect 225234 550338 225266 550894
rect 225822 550338 225854 550894
rect 225234 514894 225854 550338
rect 225234 514338 225266 514894
rect 225822 514338 225854 514894
rect 225234 478894 225854 514338
rect 225234 478338 225266 478894
rect 225822 478338 225854 478894
rect 225234 442894 225854 478338
rect 225234 442338 225266 442894
rect 225822 442338 225854 442894
rect 225234 406894 225854 442338
rect 225234 406338 225266 406894
rect 225822 406338 225854 406894
rect 225234 370894 225854 406338
rect 225234 370338 225266 370894
rect 225822 370338 225854 370894
rect 225234 334894 225854 370338
rect 225234 334338 225266 334894
rect 225822 334338 225854 334894
rect 225234 298894 225854 334338
rect 225234 298338 225266 298894
rect 225822 298338 225854 298894
rect 225234 262894 225854 298338
rect 225234 262338 225266 262894
rect 225822 262338 225854 262894
rect 225234 226894 225854 262338
rect 225234 226338 225266 226894
rect 225822 226338 225854 226894
rect 225234 190894 225854 226338
rect 225234 190338 225266 190894
rect 225822 190338 225854 190894
rect 225234 154894 225854 190338
rect 225234 154338 225266 154894
rect 225822 154338 225854 154894
rect 225234 118894 225854 154338
rect 225234 118338 225266 118894
rect 225822 118338 225854 118894
rect 225234 82894 225854 118338
rect 225234 82338 225266 82894
rect 225822 82338 225854 82894
rect 225234 46894 225854 82338
rect 225234 46338 225266 46894
rect 225822 46338 225854 46894
rect 225234 10894 225854 46338
rect 225234 10338 225266 10894
rect 225822 10338 225854 10894
rect 225234 -4186 225854 10338
rect 225234 -4742 225266 -4186
rect 225822 -4742 225854 -4186
rect 225234 -5734 225854 -4742
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711002 246986 711558
rect 247542 711002 247574 711558
rect 243234 709638 243854 709670
rect 243234 709082 243266 709638
rect 243822 709082 243854 709638
rect 239514 707718 240134 707750
rect 239514 707162 239546 707718
rect 240102 707162 240134 707718
rect 228954 698058 228986 698614
rect 229542 698058 229574 698614
rect 228954 662614 229574 698058
rect 228954 662058 228986 662614
rect 229542 662058 229574 662614
rect 228954 626614 229574 662058
rect 228954 626058 228986 626614
rect 229542 626058 229574 626614
rect 228954 590614 229574 626058
rect 228954 590058 228986 590614
rect 229542 590058 229574 590614
rect 228954 554614 229574 590058
rect 228954 554058 228986 554614
rect 229542 554058 229574 554614
rect 228954 518614 229574 554058
rect 228954 518058 228986 518614
rect 229542 518058 229574 518614
rect 228954 482614 229574 518058
rect 228954 482058 228986 482614
rect 229542 482058 229574 482614
rect 228954 446614 229574 482058
rect 228954 446058 228986 446614
rect 229542 446058 229574 446614
rect 228954 410614 229574 446058
rect 228954 410058 228986 410614
rect 229542 410058 229574 410614
rect 228954 374614 229574 410058
rect 235794 705798 236414 705830
rect 235794 705242 235826 705798
rect 236382 705242 236414 705798
rect 235794 669454 236414 705242
rect 235794 668898 235826 669454
rect 236382 668898 236414 669454
rect 235794 633454 236414 668898
rect 235794 632898 235826 633454
rect 236382 632898 236414 633454
rect 235794 597454 236414 632898
rect 235794 596898 235826 597454
rect 236382 596898 236414 597454
rect 235794 561454 236414 596898
rect 235794 560898 235826 561454
rect 236382 560898 236414 561454
rect 235794 525454 236414 560898
rect 235794 524898 235826 525454
rect 236382 524898 236414 525454
rect 235794 489454 236414 524898
rect 235794 488898 235826 489454
rect 236382 488898 236414 489454
rect 235794 453454 236414 488898
rect 235794 452898 235826 453454
rect 236382 452898 236414 453454
rect 235794 417454 236414 452898
rect 235794 416898 235826 417454
rect 236382 416898 236414 417454
rect 235794 381454 236414 416898
rect 235794 380898 235826 381454
rect 236382 380898 236414 381454
rect 235794 378000 236414 380898
rect 239514 673174 240134 707162
rect 239514 672618 239546 673174
rect 240102 672618 240134 673174
rect 239514 637174 240134 672618
rect 239514 636618 239546 637174
rect 240102 636618 240134 637174
rect 239514 601174 240134 636618
rect 239514 600618 239546 601174
rect 240102 600618 240134 601174
rect 239514 565174 240134 600618
rect 239514 564618 239546 565174
rect 240102 564618 240134 565174
rect 239514 529174 240134 564618
rect 239514 528618 239546 529174
rect 240102 528618 240134 529174
rect 239514 493174 240134 528618
rect 239514 492618 239546 493174
rect 240102 492618 240134 493174
rect 239514 457174 240134 492618
rect 239514 456618 239546 457174
rect 240102 456618 240134 457174
rect 239514 421174 240134 456618
rect 239514 420618 239546 421174
rect 240102 420618 240134 421174
rect 239514 385174 240134 420618
rect 239514 384618 239546 385174
rect 240102 384618 240134 385174
rect 239514 380000 240134 384618
rect 243234 676894 243854 709082
rect 243234 676338 243266 676894
rect 243822 676338 243854 676894
rect 243234 640894 243854 676338
rect 243234 640338 243266 640894
rect 243822 640338 243854 640894
rect 243234 604894 243854 640338
rect 243234 604338 243266 604894
rect 243822 604338 243854 604894
rect 243234 568894 243854 604338
rect 243234 568338 243266 568894
rect 243822 568338 243854 568894
rect 243234 532894 243854 568338
rect 243234 532338 243266 532894
rect 243822 532338 243854 532894
rect 243234 496894 243854 532338
rect 243234 496338 243266 496894
rect 243822 496338 243854 496894
rect 243234 460894 243854 496338
rect 243234 460338 243266 460894
rect 243822 460338 243854 460894
rect 243234 424894 243854 460338
rect 243234 424338 243266 424894
rect 243822 424338 243854 424894
rect 243234 388894 243854 424338
rect 243234 388338 243266 388894
rect 243822 388338 243854 388894
rect 243234 380000 243854 388338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710042 264986 710598
rect 265542 710042 265574 710598
rect 261234 708678 261854 709670
rect 261234 708122 261266 708678
rect 261822 708122 261854 708678
rect 257514 706758 258134 707750
rect 257514 706202 257546 706758
rect 258102 706202 258134 706758
rect 246954 680058 246986 680614
rect 247542 680058 247574 680614
rect 246954 644614 247574 680058
rect 246954 644058 246986 644614
rect 247542 644058 247574 644614
rect 246954 608614 247574 644058
rect 246954 608058 246986 608614
rect 247542 608058 247574 608614
rect 246954 572614 247574 608058
rect 246954 572058 246986 572614
rect 247542 572058 247574 572614
rect 246954 536614 247574 572058
rect 246954 536058 246986 536614
rect 247542 536058 247574 536614
rect 246954 500614 247574 536058
rect 246954 500058 246986 500614
rect 247542 500058 247574 500614
rect 246954 464614 247574 500058
rect 246954 464058 246986 464614
rect 247542 464058 247574 464614
rect 246954 428614 247574 464058
rect 246954 428058 246986 428614
rect 247542 428058 247574 428614
rect 246954 392614 247574 428058
rect 246954 392058 246986 392614
rect 247542 392058 247574 392614
rect 246954 380000 247574 392058
rect 253794 704838 254414 705830
rect 253794 704282 253826 704838
rect 254382 704282 254414 704838
rect 253794 687454 254414 704282
rect 253794 686898 253826 687454
rect 254382 686898 254414 687454
rect 253794 651454 254414 686898
rect 253794 650898 253826 651454
rect 254382 650898 254414 651454
rect 253794 615454 254414 650898
rect 253794 614898 253826 615454
rect 254382 614898 254414 615454
rect 253794 579454 254414 614898
rect 253794 578898 253826 579454
rect 254382 578898 254414 579454
rect 253794 543454 254414 578898
rect 253794 542898 253826 543454
rect 254382 542898 254414 543454
rect 253794 507454 254414 542898
rect 253794 506898 253826 507454
rect 254382 506898 254414 507454
rect 253794 471454 254414 506898
rect 253794 470898 253826 471454
rect 254382 470898 254414 471454
rect 253794 435454 254414 470898
rect 253794 434898 253826 435454
rect 254382 434898 254414 435454
rect 253794 399454 254414 434898
rect 253794 398898 253826 399454
rect 254382 398898 254414 399454
rect 253794 378000 254414 398898
rect 257514 691174 258134 706202
rect 257514 690618 257546 691174
rect 258102 690618 258134 691174
rect 257514 655174 258134 690618
rect 257514 654618 257546 655174
rect 258102 654618 258134 655174
rect 257514 619174 258134 654618
rect 257514 618618 257546 619174
rect 258102 618618 258134 619174
rect 257514 583174 258134 618618
rect 257514 582618 257546 583174
rect 258102 582618 258134 583174
rect 257514 547174 258134 582618
rect 257514 546618 257546 547174
rect 258102 546618 258134 547174
rect 257514 511174 258134 546618
rect 257514 510618 257546 511174
rect 258102 510618 258134 511174
rect 257514 475174 258134 510618
rect 257514 474618 257546 475174
rect 258102 474618 258134 475174
rect 257514 439174 258134 474618
rect 257514 438618 257546 439174
rect 258102 438618 258134 439174
rect 257514 403174 258134 438618
rect 257514 402618 257546 403174
rect 258102 402618 258134 403174
rect 257514 380000 258134 402618
rect 261234 694894 261854 708122
rect 261234 694338 261266 694894
rect 261822 694338 261854 694894
rect 261234 658894 261854 694338
rect 261234 658338 261266 658894
rect 261822 658338 261854 658894
rect 261234 622894 261854 658338
rect 261234 622338 261266 622894
rect 261822 622338 261854 622894
rect 261234 586894 261854 622338
rect 261234 586338 261266 586894
rect 261822 586338 261854 586894
rect 261234 550894 261854 586338
rect 261234 550338 261266 550894
rect 261822 550338 261854 550894
rect 261234 514894 261854 550338
rect 261234 514338 261266 514894
rect 261822 514338 261854 514894
rect 261234 478894 261854 514338
rect 261234 478338 261266 478894
rect 261822 478338 261854 478894
rect 261234 442894 261854 478338
rect 261234 442338 261266 442894
rect 261822 442338 261854 442894
rect 261234 406894 261854 442338
rect 261234 406338 261266 406894
rect 261822 406338 261854 406894
rect 261234 380000 261854 406338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711002 282986 711558
rect 283542 711002 283574 711558
rect 279234 709638 279854 709670
rect 279234 709082 279266 709638
rect 279822 709082 279854 709638
rect 275514 707718 276134 707750
rect 275514 707162 275546 707718
rect 276102 707162 276134 707718
rect 264954 698058 264986 698614
rect 265542 698058 265574 698614
rect 264954 662614 265574 698058
rect 264954 662058 264986 662614
rect 265542 662058 265574 662614
rect 264954 626614 265574 662058
rect 264954 626058 264986 626614
rect 265542 626058 265574 626614
rect 264954 590614 265574 626058
rect 264954 590058 264986 590614
rect 265542 590058 265574 590614
rect 264954 554614 265574 590058
rect 264954 554058 264986 554614
rect 265542 554058 265574 554614
rect 264954 518614 265574 554058
rect 264954 518058 264986 518614
rect 265542 518058 265574 518614
rect 264954 482614 265574 518058
rect 264954 482058 264986 482614
rect 265542 482058 265574 482614
rect 264954 446614 265574 482058
rect 264954 446058 264986 446614
rect 265542 446058 265574 446614
rect 264954 410614 265574 446058
rect 264954 410058 264986 410614
rect 265542 410058 265574 410614
rect 264954 380000 265574 410058
rect 271794 705798 272414 705830
rect 271794 705242 271826 705798
rect 272382 705242 272414 705798
rect 271794 669454 272414 705242
rect 271794 668898 271826 669454
rect 272382 668898 272414 669454
rect 271794 633454 272414 668898
rect 271794 632898 271826 633454
rect 272382 632898 272414 633454
rect 271794 597454 272414 632898
rect 271794 596898 271826 597454
rect 272382 596898 272414 597454
rect 271794 561454 272414 596898
rect 271794 560898 271826 561454
rect 272382 560898 272414 561454
rect 271794 525454 272414 560898
rect 271794 524898 271826 525454
rect 272382 524898 272414 525454
rect 271794 489454 272414 524898
rect 271794 488898 271826 489454
rect 272382 488898 272414 489454
rect 271794 453454 272414 488898
rect 271794 452898 271826 453454
rect 272382 452898 272414 453454
rect 271794 417454 272414 452898
rect 271794 416898 271826 417454
rect 272382 416898 272414 417454
rect 271794 381454 272414 416898
rect 271794 380898 271826 381454
rect 272382 380898 272414 381454
rect 271794 378000 272414 380898
rect 275514 673174 276134 707162
rect 275514 672618 275546 673174
rect 276102 672618 276134 673174
rect 275514 637174 276134 672618
rect 275514 636618 275546 637174
rect 276102 636618 276134 637174
rect 275514 601174 276134 636618
rect 275514 600618 275546 601174
rect 276102 600618 276134 601174
rect 275514 565174 276134 600618
rect 275514 564618 275546 565174
rect 276102 564618 276134 565174
rect 275514 529174 276134 564618
rect 275514 528618 275546 529174
rect 276102 528618 276134 529174
rect 275514 493174 276134 528618
rect 275514 492618 275546 493174
rect 276102 492618 276134 493174
rect 275514 457174 276134 492618
rect 275514 456618 275546 457174
rect 276102 456618 276134 457174
rect 275514 421174 276134 456618
rect 275514 420618 275546 421174
rect 276102 420618 276134 421174
rect 275514 385174 276134 420618
rect 275514 384618 275546 385174
rect 276102 384618 276134 385174
rect 275514 380000 276134 384618
rect 279234 676894 279854 709082
rect 279234 676338 279266 676894
rect 279822 676338 279854 676894
rect 279234 640894 279854 676338
rect 279234 640338 279266 640894
rect 279822 640338 279854 640894
rect 279234 604894 279854 640338
rect 279234 604338 279266 604894
rect 279822 604338 279854 604894
rect 279234 568894 279854 604338
rect 279234 568338 279266 568894
rect 279822 568338 279854 568894
rect 279234 532894 279854 568338
rect 279234 532338 279266 532894
rect 279822 532338 279854 532894
rect 279234 496894 279854 532338
rect 279234 496338 279266 496894
rect 279822 496338 279854 496894
rect 279234 460894 279854 496338
rect 279234 460338 279266 460894
rect 279822 460338 279854 460894
rect 279234 424894 279854 460338
rect 279234 424338 279266 424894
rect 279822 424338 279854 424894
rect 279234 388894 279854 424338
rect 279234 388338 279266 388894
rect 279822 388338 279854 388894
rect 279234 380000 279854 388338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710042 300986 710598
rect 301542 710042 301574 710598
rect 297234 708678 297854 709670
rect 297234 708122 297266 708678
rect 297822 708122 297854 708678
rect 293514 706758 294134 707750
rect 293514 706202 293546 706758
rect 294102 706202 294134 706758
rect 282954 680058 282986 680614
rect 283542 680058 283574 680614
rect 282954 644614 283574 680058
rect 282954 644058 282986 644614
rect 283542 644058 283574 644614
rect 282954 608614 283574 644058
rect 282954 608058 282986 608614
rect 283542 608058 283574 608614
rect 282954 572614 283574 608058
rect 282954 572058 282986 572614
rect 283542 572058 283574 572614
rect 282954 536614 283574 572058
rect 282954 536058 282986 536614
rect 283542 536058 283574 536614
rect 282954 500614 283574 536058
rect 282954 500058 282986 500614
rect 283542 500058 283574 500614
rect 282954 464614 283574 500058
rect 282954 464058 282986 464614
rect 283542 464058 283574 464614
rect 282954 428614 283574 464058
rect 282954 428058 282986 428614
rect 283542 428058 283574 428614
rect 282954 392614 283574 428058
rect 282954 392058 282986 392614
rect 283542 392058 283574 392614
rect 282954 380000 283574 392058
rect 289794 704838 290414 705830
rect 289794 704282 289826 704838
rect 290382 704282 290414 704838
rect 289794 687454 290414 704282
rect 289794 686898 289826 687454
rect 290382 686898 290414 687454
rect 289794 651454 290414 686898
rect 289794 650898 289826 651454
rect 290382 650898 290414 651454
rect 289794 615454 290414 650898
rect 289794 614898 289826 615454
rect 290382 614898 290414 615454
rect 289794 579454 290414 614898
rect 289794 578898 289826 579454
rect 290382 578898 290414 579454
rect 289794 543454 290414 578898
rect 289794 542898 289826 543454
rect 290382 542898 290414 543454
rect 289794 507454 290414 542898
rect 289794 506898 289826 507454
rect 290382 506898 290414 507454
rect 289794 471454 290414 506898
rect 289794 470898 289826 471454
rect 290382 470898 290414 471454
rect 289794 435454 290414 470898
rect 289794 434898 289826 435454
rect 290382 434898 290414 435454
rect 289794 399454 290414 434898
rect 289794 398898 289826 399454
rect 290382 398898 290414 399454
rect 289794 378000 290414 398898
rect 293514 691174 294134 706202
rect 293514 690618 293546 691174
rect 294102 690618 294134 691174
rect 293514 655174 294134 690618
rect 293514 654618 293546 655174
rect 294102 654618 294134 655174
rect 293514 619174 294134 654618
rect 293514 618618 293546 619174
rect 294102 618618 294134 619174
rect 293514 583174 294134 618618
rect 293514 582618 293546 583174
rect 294102 582618 294134 583174
rect 293514 547174 294134 582618
rect 293514 546618 293546 547174
rect 294102 546618 294134 547174
rect 293514 511174 294134 546618
rect 293514 510618 293546 511174
rect 294102 510618 294134 511174
rect 293514 475174 294134 510618
rect 293514 474618 293546 475174
rect 294102 474618 294134 475174
rect 293514 439174 294134 474618
rect 293514 438618 293546 439174
rect 294102 438618 294134 439174
rect 293514 403174 294134 438618
rect 293514 402618 293546 403174
rect 294102 402618 294134 403174
rect 293514 380000 294134 402618
rect 297234 694894 297854 708122
rect 297234 694338 297266 694894
rect 297822 694338 297854 694894
rect 297234 658894 297854 694338
rect 297234 658338 297266 658894
rect 297822 658338 297854 658894
rect 297234 622894 297854 658338
rect 297234 622338 297266 622894
rect 297822 622338 297854 622894
rect 297234 586894 297854 622338
rect 297234 586338 297266 586894
rect 297822 586338 297854 586894
rect 297234 550894 297854 586338
rect 297234 550338 297266 550894
rect 297822 550338 297854 550894
rect 297234 514894 297854 550338
rect 297234 514338 297266 514894
rect 297822 514338 297854 514894
rect 297234 478894 297854 514338
rect 297234 478338 297266 478894
rect 297822 478338 297854 478894
rect 297234 442894 297854 478338
rect 297234 442338 297266 442894
rect 297822 442338 297854 442894
rect 297234 406894 297854 442338
rect 297234 406338 297266 406894
rect 297822 406338 297854 406894
rect 237235 377364 237301 377365
rect 237235 377300 237236 377364
rect 237300 377300 237301 377364
rect 237235 377299 237301 377300
rect 238523 377364 238589 377365
rect 238523 377300 238524 377364
rect 238588 377300 238589 377364
rect 238523 377299 238589 377300
rect 241283 377364 241349 377365
rect 241283 377300 241284 377364
rect 241348 377300 241349 377364
rect 241283 377299 241349 377300
rect 242755 377364 242821 377365
rect 242755 377300 242756 377364
rect 242820 377300 242821 377364
rect 242755 377299 242821 377300
rect 244043 377364 244109 377365
rect 244043 377300 244044 377364
rect 244108 377300 244109 377364
rect 244043 377299 244109 377300
rect 285811 377364 285877 377365
rect 285811 377300 285812 377364
rect 285876 377300 285877 377364
rect 285811 377299 285877 377300
rect 287099 377364 287165 377365
rect 287099 377300 287100 377364
rect 287164 377300 287165 377364
rect 287099 377299 287165 377300
rect 288387 377364 288453 377365
rect 288387 377300 288388 377364
rect 288452 377300 288453 377364
rect 288387 377299 288453 377300
rect 290595 377364 290661 377365
rect 290595 377300 290596 377364
rect 290660 377300 290661 377364
rect 290595 377299 290661 377300
rect 291147 377364 291213 377365
rect 291147 377300 291148 377364
rect 291212 377300 291213 377364
rect 291147 377299 291213 377300
rect 292619 377364 292685 377365
rect 292619 377300 292620 377364
rect 292684 377300 292685 377364
rect 292619 377299 292685 377300
rect 228954 374058 228986 374614
rect 229542 374058 229574 374614
rect 228954 338614 229574 374058
rect 228954 338058 228986 338614
rect 229542 338058 229574 338614
rect 228954 302614 229574 338058
rect 228954 302058 228986 302614
rect 229542 302058 229574 302614
rect 228954 266614 229574 302058
rect 228954 266058 228986 266614
rect 229542 266058 229574 266614
rect 228954 230614 229574 266058
rect 228954 230058 228986 230614
rect 229542 230058 229574 230614
rect 228954 194614 229574 230058
rect 228954 194058 228986 194614
rect 229542 194058 229574 194614
rect 228954 158614 229574 194058
rect 228954 158058 228986 158614
rect 229542 158058 229574 158614
rect 228954 122614 229574 158058
rect 228954 122058 228986 122614
rect 229542 122058 229574 122614
rect 228954 86614 229574 122058
rect 228954 86058 228986 86614
rect 229542 86058 229574 86614
rect 228954 50614 229574 86058
rect 228954 50058 228986 50614
rect 229542 50058 229574 50614
rect 228954 14614 229574 50058
rect 228954 14058 228986 14614
rect 229542 14058 229574 14614
rect 210954 -7622 210986 -7066
rect 211542 -7622 211574 -7066
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 309454 236414 338000
rect 235794 308898 235826 309454
rect 236382 308898 236414 309454
rect 235794 273454 236414 308898
rect 235794 272898 235826 273454
rect 236382 272898 236414 273454
rect 235794 237454 236414 272898
rect 235794 236898 235826 237454
rect 236382 236898 236414 237454
rect 235794 201454 236414 236898
rect 235794 200898 235826 201454
rect 236382 200898 236414 201454
rect 235794 165454 236414 200898
rect 235794 164898 235826 165454
rect 236382 164898 236414 165454
rect 235794 129454 236414 164898
rect 235794 128898 235826 129454
rect 236382 128898 236414 129454
rect 235794 93454 236414 128898
rect 235794 92898 235826 93454
rect 236382 92898 236414 93454
rect 235794 57454 236414 92898
rect 235794 56898 235826 57454
rect 236382 56898 236414 57454
rect 235794 21454 236414 56898
rect 235794 20898 235826 21454
rect 236382 20898 236414 21454
rect 235794 -1306 236414 20898
rect 237238 19413 237298 377299
rect 238526 59397 238586 377299
rect 239208 363454 239528 363486
rect 239208 363218 239250 363454
rect 239486 363218 239528 363454
rect 239208 363134 239528 363218
rect 239208 362898 239250 363134
rect 239486 362898 239528 363134
rect 239208 362866 239528 362898
rect 239514 313174 240134 336000
rect 239514 312618 239546 313174
rect 240102 312618 240134 313174
rect 239514 277174 240134 312618
rect 239514 276618 239546 277174
rect 240102 276618 240134 277174
rect 239514 241174 240134 276618
rect 239514 240618 239546 241174
rect 240102 240618 240134 241174
rect 239514 205174 240134 240618
rect 239514 204618 239546 205174
rect 240102 204618 240134 205174
rect 239514 169174 240134 204618
rect 239514 168618 239546 169174
rect 240102 168618 240134 169174
rect 239514 133174 240134 168618
rect 241286 138141 241346 377299
rect 242758 178125 242818 377299
rect 243234 316894 243854 336000
rect 243234 316338 243266 316894
rect 243822 316338 243854 316894
rect 243234 280894 243854 316338
rect 243234 280338 243266 280894
rect 243822 280338 243854 280894
rect 243234 244894 243854 280338
rect 243234 244338 243266 244894
rect 243822 244338 243854 244894
rect 243234 208894 243854 244338
rect 244046 218109 244106 377299
rect 269928 363454 270248 363486
rect 269928 363218 269970 363454
rect 270206 363218 270248 363454
rect 269928 363134 270248 363218
rect 269928 362898 269970 363134
rect 270206 362898 270248 363134
rect 269928 362866 270248 362898
rect 254568 345454 254888 345486
rect 254568 345218 254610 345454
rect 254846 345218 254888 345454
rect 254568 345134 254888 345218
rect 254568 344898 254610 345134
rect 254846 344898 254888 345134
rect 254568 344866 254888 344898
rect 285288 345454 285608 345486
rect 285288 345218 285330 345454
rect 285566 345218 285608 345454
rect 285288 345134 285608 345218
rect 285288 344898 285330 345134
rect 285566 344898 285608 345134
rect 285288 344866 285608 344898
rect 246954 320614 247574 336000
rect 246954 320058 246986 320614
rect 247542 320058 247574 320614
rect 246954 284614 247574 320058
rect 246954 284058 246986 284614
rect 247542 284058 247574 284614
rect 246954 248614 247574 284058
rect 246954 248058 246986 248614
rect 247542 248058 247574 248614
rect 244043 218108 244109 218109
rect 244043 218044 244044 218108
rect 244108 218044 244109 218108
rect 244043 218043 244109 218044
rect 243234 208338 243266 208894
rect 243822 208338 243854 208894
rect 242755 178124 242821 178125
rect 242755 178060 242756 178124
rect 242820 178060 242821 178124
rect 242755 178059 242821 178060
rect 243234 172894 243854 208338
rect 243234 172338 243266 172894
rect 243822 172338 243854 172894
rect 241283 138140 241349 138141
rect 241283 138076 241284 138140
rect 241348 138076 241349 138140
rect 241283 138075 241349 138076
rect 239514 132618 239546 133174
rect 240102 132618 240134 133174
rect 239514 97174 240134 132618
rect 239514 96618 239546 97174
rect 240102 96618 240134 97174
rect 239514 61174 240134 96618
rect 239514 60618 239546 61174
rect 240102 60618 240134 61174
rect 238523 59396 238589 59397
rect 238523 59332 238524 59396
rect 238588 59332 238589 59396
rect 238523 59331 238589 59332
rect 239514 25174 240134 60618
rect 239514 24618 239546 25174
rect 240102 24618 240134 25174
rect 237235 19412 237301 19413
rect 237235 19348 237236 19412
rect 237300 19348 237301 19412
rect 237235 19347 237301 19348
rect 235794 -1862 235826 -1306
rect 236382 -1862 236414 -1306
rect 235794 -1894 236414 -1862
rect 239514 -3226 240134 24618
rect 239514 -3782 239546 -3226
rect 240102 -3782 240134 -3226
rect 239514 -3814 240134 -3782
rect 243234 136894 243854 172338
rect 243234 136338 243266 136894
rect 243822 136338 243854 136894
rect 243234 100894 243854 136338
rect 243234 100338 243266 100894
rect 243822 100338 243854 100894
rect 243234 64894 243854 100338
rect 243234 64338 243266 64894
rect 243822 64338 243854 64894
rect 243234 28894 243854 64338
rect 243234 28338 243266 28894
rect 243822 28338 243854 28894
rect 243234 -5146 243854 28338
rect 243234 -5702 243266 -5146
rect 243822 -5702 243854 -5146
rect 243234 -5734 243854 -5702
rect 246954 212614 247574 248058
rect 246954 212058 246986 212614
rect 247542 212058 247574 212614
rect 246954 176614 247574 212058
rect 246954 176058 246986 176614
rect 247542 176058 247574 176614
rect 246954 140614 247574 176058
rect 246954 140058 246986 140614
rect 247542 140058 247574 140614
rect 246954 104614 247574 140058
rect 246954 104058 246986 104614
rect 247542 104058 247574 104614
rect 246954 68614 247574 104058
rect 246954 68058 246986 68614
rect 247542 68058 247574 68614
rect 246954 32614 247574 68058
rect 246954 32058 246986 32614
rect 247542 32058 247574 32614
rect 228954 -6662 228986 -6106
rect 229542 -6662 229574 -6106
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 327454 254414 338000
rect 253794 326898 253826 327454
rect 254382 326898 254414 327454
rect 253794 291454 254414 326898
rect 253794 290898 253826 291454
rect 254382 290898 254414 291454
rect 253794 255454 254414 290898
rect 253794 254898 253826 255454
rect 254382 254898 254414 255454
rect 253794 219454 254414 254898
rect 253794 218898 253826 219454
rect 254382 218898 254414 219454
rect 253794 183454 254414 218898
rect 253794 182898 253826 183454
rect 254382 182898 254414 183454
rect 253794 147454 254414 182898
rect 253794 146898 253826 147454
rect 254382 146898 254414 147454
rect 253794 111454 254414 146898
rect 253794 110898 253826 111454
rect 254382 110898 254414 111454
rect 253794 75454 254414 110898
rect 253794 74898 253826 75454
rect 254382 74898 254414 75454
rect 253794 39454 254414 74898
rect 253794 38898 253826 39454
rect 254382 38898 254414 39454
rect 253794 3454 254414 38898
rect 253794 2898 253826 3454
rect 254382 2898 254414 3454
rect 253794 -346 254414 2898
rect 253794 -902 253826 -346
rect 254382 -902 254414 -346
rect 253794 -1894 254414 -902
rect 257514 331174 258134 336000
rect 257514 330618 257546 331174
rect 258102 330618 258134 331174
rect 257514 295174 258134 330618
rect 257514 294618 257546 295174
rect 258102 294618 258134 295174
rect 257514 259174 258134 294618
rect 257514 258618 257546 259174
rect 258102 258618 258134 259174
rect 257514 223174 258134 258618
rect 257514 222618 257546 223174
rect 258102 222618 258134 223174
rect 257514 187174 258134 222618
rect 257514 186618 257546 187174
rect 258102 186618 258134 187174
rect 257514 151174 258134 186618
rect 257514 150618 257546 151174
rect 258102 150618 258134 151174
rect 257514 115174 258134 150618
rect 257514 114618 257546 115174
rect 258102 114618 258134 115174
rect 257514 79174 258134 114618
rect 257514 78618 257546 79174
rect 258102 78618 258134 79174
rect 257514 43174 258134 78618
rect 257514 42618 257546 43174
rect 258102 42618 258134 43174
rect 257514 7174 258134 42618
rect 257514 6618 257546 7174
rect 258102 6618 258134 7174
rect 257514 -2266 258134 6618
rect 257514 -2822 257546 -2266
rect 258102 -2822 258134 -2266
rect 257514 -3814 258134 -2822
rect 261234 334894 261854 336000
rect 261234 334338 261266 334894
rect 261822 334338 261854 334894
rect 261234 298894 261854 334338
rect 261234 298338 261266 298894
rect 261822 298338 261854 298894
rect 261234 262894 261854 298338
rect 261234 262338 261266 262894
rect 261822 262338 261854 262894
rect 261234 226894 261854 262338
rect 261234 226338 261266 226894
rect 261822 226338 261854 226894
rect 261234 190894 261854 226338
rect 261234 190338 261266 190894
rect 261822 190338 261854 190894
rect 261234 154894 261854 190338
rect 261234 154338 261266 154894
rect 261822 154338 261854 154894
rect 261234 118894 261854 154338
rect 261234 118338 261266 118894
rect 261822 118338 261854 118894
rect 261234 82894 261854 118338
rect 261234 82338 261266 82894
rect 261822 82338 261854 82894
rect 261234 46894 261854 82338
rect 261234 46338 261266 46894
rect 261822 46338 261854 46894
rect 261234 10894 261854 46338
rect 261234 10338 261266 10894
rect 261822 10338 261854 10894
rect 261234 -4186 261854 10338
rect 261234 -4742 261266 -4186
rect 261822 -4742 261854 -4186
rect 261234 -5734 261854 -4742
rect 264954 302614 265574 336000
rect 264954 302058 264986 302614
rect 265542 302058 265574 302614
rect 264954 266614 265574 302058
rect 264954 266058 264986 266614
rect 265542 266058 265574 266614
rect 264954 230614 265574 266058
rect 264954 230058 264986 230614
rect 265542 230058 265574 230614
rect 264954 194614 265574 230058
rect 264954 194058 264986 194614
rect 265542 194058 265574 194614
rect 264954 158614 265574 194058
rect 264954 158058 264986 158614
rect 265542 158058 265574 158614
rect 264954 122614 265574 158058
rect 264954 122058 264986 122614
rect 265542 122058 265574 122614
rect 264954 86614 265574 122058
rect 264954 86058 264986 86614
rect 265542 86058 265574 86614
rect 264954 50614 265574 86058
rect 264954 50058 264986 50614
rect 265542 50058 265574 50614
rect 264954 14614 265574 50058
rect 264954 14058 264986 14614
rect 265542 14058 265574 14614
rect 246954 -7622 246986 -7066
rect 247542 -7622 247574 -7066
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 309454 272414 338000
rect 271794 308898 271826 309454
rect 272382 308898 272414 309454
rect 271794 273454 272414 308898
rect 271794 272898 271826 273454
rect 272382 272898 272414 273454
rect 271794 237454 272414 272898
rect 271794 236898 271826 237454
rect 272382 236898 272414 237454
rect 271794 201454 272414 236898
rect 271794 200898 271826 201454
rect 272382 200898 272414 201454
rect 271794 165454 272414 200898
rect 271794 164898 271826 165454
rect 272382 164898 272414 165454
rect 271794 129454 272414 164898
rect 271794 128898 271826 129454
rect 272382 128898 272414 129454
rect 271794 93454 272414 128898
rect 271794 92898 271826 93454
rect 272382 92898 272414 93454
rect 271794 57454 272414 92898
rect 271794 56898 271826 57454
rect 272382 56898 272414 57454
rect 271794 21454 272414 56898
rect 271794 20898 271826 21454
rect 272382 20898 272414 21454
rect 271794 -1306 272414 20898
rect 271794 -1862 271826 -1306
rect 272382 -1862 272414 -1306
rect 271794 -1894 272414 -1862
rect 275514 313174 276134 336000
rect 275514 312618 275546 313174
rect 276102 312618 276134 313174
rect 275514 277174 276134 312618
rect 275514 276618 275546 277174
rect 276102 276618 276134 277174
rect 275514 241174 276134 276618
rect 275514 240618 275546 241174
rect 276102 240618 276134 241174
rect 275514 205174 276134 240618
rect 275514 204618 275546 205174
rect 276102 204618 276134 205174
rect 275514 169174 276134 204618
rect 275514 168618 275546 169174
rect 276102 168618 276134 169174
rect 275514 133174 276134 168618
rect 275514 132618 275546 133174
rect 276102 132618 276134 133174
rect 275514 97174 276134 132618
rect 275514 96618 275546 97174
rect 276102 96618 276134 97174
rect 275514 61174 276134 96618
rect 275514 60618 275546 61174
rect 276102 60618 276134 61174
rect 275514 25174 276134 60618
rect 275514 24618 275546 25174
rect 276102 24618 276134 25174
rect 275514 -3226 276134 24618
rect 275514 -3782 275546 -3226
rect 276102 -3782 276134 -3226
rect 275514 -3814 276134 -3782
rect 279234 316894 279854 336000
rect 279234 316338 279266 316894
rect 279822 316338 279854 316894
rect 279234 280894 279854 316338
rect 279234 280338 279266 280894
rect 279822 280338 279854 280894
rect 279234 244894 279854 280338
rect 279234 244338 279266 244894
rect 279822 244338 279854 244894
rect 279234 208894 279854 244338
rect 279234 208338 279266 208894
rect 279822 208338 279854 208894
rect 279234 172894 279854 208338
rect 279234 172338 279266 172894
rect 279822 172338 279854 172894
rect 279234 136894 279854 172338
rect 279234 136338 279266 136894
rect 279822 136338 279854 136894
rect 279234 100894 279854 136338
rect 279234 100338 279266 100894
rect 279822 100338 279854 100894
rect 279234 64894 279854 100338
rect 279234 64338 279266 64894
rect 279822 64338 279854 64894
rect 279234 28894 279854 64338
rect 279234 28338 279266 28894
rect 279822 28338 279854 28894
rect 279234 -5146 279854 28338
rect 279234 -5702 279266 -5146
rect 279822 -5702 279854 -5146
rect 279234 -5734 279854 -5702
rect 282954 320614 283574 336000
rect 282954 320058 282986 320614
rect 283542 320058 283574 320614
rect 282954 284614 283574 320058
rect 282954 284058 282986 284614
rect 283542 284058 283574 284614
rect 282954 248614 283574 284058
rect 285814 255237 285874 377299
rect 285811 255236 285877 255237
rect 285811 255172 285812 255236
rect 285876 255172 285877 255236
rect 285811 255171 285877 255172
rect 282954 248058 282986 248614
rect 283542 248058 283574 248614
rect 282954 212614 283574 248058
rect 282954 212058 282986 212614
rect 283542 212058 283574 212614
rect 282954 176614 283574 212058
rect 287102 202877 287162 377299
rect 287099 202876 287165 202877
rect 287099 202812 287100 202876
rect 287164 202812 287165 202876
rect 287099 202811 287165 202812
rect 282954 176058 282986 176614
rect 283542 176058 283574 176614
rect 282954 140614 283574 176058
rect 282954 140058 282986 140614
rect 283542 140058 283574 140614
rect 282954 104614 283574 140058
rect 288390 138005 288450 377299
rect 289794 327454 290414 338000
rect 289794 326898 289826 327454
rect 290382 326898 290414 327454
rect 289794 291454 290414 326898
rect 289794 290898 289826 291454
rect 290382 290898 290414 291454
rect 289794 255454 290414 290898
rect 289794 254898 289826 255454
rect 290382 254898 290414 255454
rect 289794 219454 290414 254898
rect 289794 218898 289826 219454
rect 290382 218898 290414 219454
rect 289794 183454 290414 218898
rect 289794 182898 289826 183454
rect 290382 182898 290414 183454
rect 289794 147454 290414 182898
rect 290598 150381 290658 377299
rect 290595 150380 290661 150381
rect 290595 150316 290596 150380
rect 290660 150316 290661 150380
rect 290595 150315 290661 150316
rect 289794 146898 289826 147454
rect 290382 146898 290414 147454
rect 288387 138004 288453 138005
rect 288387 137940 288388 138004
rect 288452 137940 288453 138004
rect 288387 137939 288453 137940
rect 282954 104058 282986 104614
rect 283542 104058 283574 104614
rect 282954 68614 283574 104058
rect 282954 68058 282986 68614
rect 283542 68058 283574 68614
rect 282954 32614 283574 68058
rect 282954 32058 282986 32614
rect 283542 32058 283574 32614
rect 264954 -6662 264986 -6106
rect 265542 -6662 265574 -6106
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 111454 290414 146898
rect 289794 110898 289826 111454
rect 290382 110898 290414 111454
rect 289794 75454 290414 110898
rect 291150 97885 291210 377299
rect 291147 97884 291213 97885
rect 291147 97820 291148 97884
rect 291212 97820 291213 97884
rect 291147 97819 291213 97820
rect 289794 74898 289826 75454
rect 290382 74898 290414 75454
rect 289794 39454 290414 74898
rect 292622 59261 292682 377299
rect 297234 370894 297854 406338
rect 297234 370338 297266 370894
rect 297822 370338 297854 370894
rect 293514 331174 294134 336000
rect 293514 330618 293546 331174
rect 294102 330618 294134 331174
rect 293514 295174 294134 330618
rect 293514 294618 293546 295174
rect 294102 294618 294134 295174
rect 293514 259174 294134 294618
rect 293514 258618 293546 259174
rect 294102 258618 294134 259174
rect 293514 223174 294134 258618
rect 293514 222618 293546 223174
rect 294102 222618 294134 223174
rect 293514 187174 294134 222618
rect 293514 186618 293546 187174
rect 294102 186618 294134 187174
rect 293514 151174 294134 186618
rect 293514 150618 293546 151174
rect 294102 150618 294134 151174
rect 293514 115174 294134 150618
rect 293514 114618 293546 115174
rect 294102 114618 294134 115174
rect 293514 79174 294134 114618
rect 293514 78618 293546 79174
rect 294102 78618 294134 79174
rect 292619 59260 292685 59261
rect 292619 59196 292620 59260
rect 292684 59196 292685 59260
rect 292619 59195 292685 59196
rect 289794 38898 289826 39454
rect 290382 38898 290414 39454
rect 289794 3454 290414 38898
rect 289794 2898 289826 3454
rect 290382 2898 290414 3454
rect 289794 -346 290414 2898
rect 289794 -902 289826 -346
rect 290382 -902 290414 -346
rect 289794 -1894 290414 -902
rect 293514 43174 294134 78618
rect 293514 42618 293546 43174
rect 294102 42618 294134 43174
rect 293514 7174 294134 42618
rect 293514 6618 293546 7174
rect 294102 6618 294134 7174
rect 293514 -2266 294134 6618
rect 293514 -2822 293546 -2266
rect 294102 -2822 294134 -2266
rect 293514 -3814 294134 -2822
rect 297234 334894 297854 370338
rect 297234 334338 297266 334894
rect 297822 334338 297854 334894
rect 297234 298894 297854 334338
rect 297234 298338 297266 298894
rect 297822 298338 297854 298894
rect 297234 262894 297854 298338
rect 297234 262338 297266 262894
rect 297822 262338 297854 262894
rect 297234 226894 297854 262338
rect 297234 226338 297266 226894
rect 297822 226338 297854 226894
rect 297234 190894 297854 226338
rect 297234 190338 297266 190894
rect 297822 190338 297854 190894
rect 297234 154894 297854 190338
rect 297234 154338 297266 154894
rect 297822 154338 297854 154894
rect 297234 118894 297854 154338
rect 297234 118338 297266 118894
rect 297822 118338 297854 118894
rect 297234 82894 297854 118338
rect 297234 82338 297266 82894
rect 297822 82338 297854 82894
rect 297234 46894 297854 82338
rect 297234 46338 297266 46894
rect 297822 46338 297854 46894
rect 297234 10894 297854 46338
rect 297234 10338 297266 10894
rect 297822 10338 297854 10894
rect 297234 -4186 297854 10338
rect 297234 -4742 297266 -4186
rect 297822 -4742 297854 -4186
rect 297234 -5734 297854 -4742
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711002 318986 711558
rect 319542 711002 319574 711558
rect 315234 709638 315854 709670
rect 315234 709082 315266 709638
rect 315822 709082 315854 709638
rect 311514 707718 312134 707750
rect 311514 707162 311546 707718
rect 312102 707162 312134 707718
rect 300954 698058 300986 698614
rect 301542 698058 301574 698614
rect 300954 662614 301574 698058
rect 300954 662058 300986 662614
rect 301542 662058 301574 662614
rect 300954 626614 301574 662058
rect 300954 626058 300986 626614
rect 301542 626058 301574 626614
rect 300954 590614 301574 626058
rect 300954 590058 300986 590614
rect 301542 590058 301574 590614
rect 300954 554614 301574 590058
rect 300954 554058 300986 554614
rect 301542 554058 301574 554614
rect 300954 518614 301574 554058
rect 300954 518058 300986 518614
rect 301542 518058 301574 518614
rect 300954 482614 301574 518058
rect 300954 482058 300986 482614
rect 301542 482058 301574 482614
rect 300954 446614 301574 482058
rect 300954 446058 300986 446614
rect 301542 446058 301574 446614
rect 300954 410614 301574 446058
rect 300954 410058 300986 410614
rect 301542 410058 301574 410614
rect 300954 374614 301574 410058
rect 300954 374058 300986 374614
rect 301542 374058 301574 374614
rect 300954 338614 301574 374058
rect 300954 338058 300986 338614
rect 301542 338058 301574 338614
rect 300954 302614 301574 338058
rect 300954 302058 300986 302614
rect 301542 302058 301574 302614
rect 300954 266614 301574 302058
rect 300954 266058 300986 266614
rect 301542 266058 301574 266614
rect 300954 230614 301574 266058
rect 300954 230058 300986 230614
rect 301542 230058 301574 230614
rect 300954 194614 301574 230058
rect 300954 194058 300986 194614
rect 301542 194058 301574 194614
rect 300954 158614 301574 194058
rect 300954 158058 300986 158614
rect 301542 158058 301574 158614
rect 300954 122614 301574 158058
rect 300954 122058 300986 122614
rect 301542 122058 301574 122614
rect 300954 86614 301574 122058
rect 300954 86058 300986 86614
rect 301542 86058 301574 86614
rect 300954 50614 301574 86058
rect 300954 50058 300986 50614
rect 301542 50058 301574 50614
rect 300954 14614 301574 50058
rect 300954 14058 300986 14614
rect 301542 14058 301574 14614
rect 282954 -7622 282986 -7066
rect 283542 -7622 283574 -7066
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 705798 308414 705830
rect 307794 705242 307826 705798
rect 308382 705242 308414 705798
rect 307794 669454 308414 705242
rect 307794 668898 307826 669454
rect 308382 668898 308414 669454
rect 307794 633454 308414 668898
rect 307794 632898 307826 633454
rect 308382 632898 308414 633454
rect 307794 597454 308414 632898
rect 307794 596898 307826 597454
rect 308382 596898 308414 597454
rect 307794 561454 308414 596898
rect 307794 560898 307826 561454
rect 308382 560898 308414 561454
rect 307794 525454 308414 560898
rect 307794 524898 307826 525454
rect 308382 524898 308414 525454
rect 307794 489454 308414 524898
rect 307794 488898 307826 489454
rect 308382 488898 308414 489454
rect 307794 453454 308414 488898
rect 307794 452898 307826 453454
rect 308382 452898 308414 453454
rect 307794 417454 308414 452898
rect 307794 416898 307826 417454
rect 308382 416898 308414 417454
rect 307794 381454 308414 416898
rect 307794 380898 307826 381454
rect 308382 380898 308414 381454
rect 307794 345454 308414 380898
rect 307794 344898 307826 345454
rect 308382 344898 308414 345454
rect 307794 309454 308414 344898
rect 307794 308898 307826 309454
rect 308382 308898 308414 309454
rect 307794 273454 308414 308898
rect 307794 272898 307826 273454
rect 308382 272898 308414 273454
rect 307794 237454 308414 272898
rect 307794 236898 307826 237454
rect 308382 236898 308414 237454
rect 307794 201454 308414 236898
rect 307794 200898 307826 201454
rect 308382 200898 308414 201454
rect 307794 165454 308414 200898
rect 307794 164898 307826 165454
rect 308382 164898 308414 165454
rect 307794 129454 308414 164898
rect 307794 128898 307826 129454
rect 308382 128898 308414 129454
rect 307794 93454 308414 128898
rect 307794 92898 307826 93454
rect 308382 92898 308414 93454
rect 307794 57454 308414 92898
rect 307794 56898 307826 57454
rect 308382 56898 308414 57454
rect 307794 21454 308414 56898
rect 307794 20898 307826 21454
rect 308382 20898 308414 21454
rect 307794 -1306 308414 20898
rect 307794 -1862 307826 -1306
rect 308382 -1862 308414 -1306
rect 307794 -1894 308414 -1862
rect 311514 673174 312134 707162
rect 311514 672618 311546 673174
rect 312102 672618 312134 673174
rect 311514 637174 312134 672618
rect 311514 636618 311546 637174
rect 312102 636618 312134 637174
rect 311514 601174 312134 636618
rect 311514 600618 311546 601174
rect 312102 600618 312134 601174
rect 311514 565174 312134 600618
rect 311514 564618 311546 565174
rect 312102 564618 312134 565174
rect 311514 529174 312134 564618
rect 311514 528618 311546 529174
rect 312102 528618 312134 529174
rect 311514 493174 312134 528618
rect 311514 492618 311546 493174
rect 312102 492618 312134 493174
rect 311514 457174 312134 492618
rect 311514 456618 311546 457174
rect 312102 456618 312134 457174
rect 311514 421174 312134 456618
rect 311514 420618 311546 421174
rect 312102 420618 312134 421174
rect 311514 385174 312134 420618
rect 311514 384618 311546 385174
rect 312102 384618 312134 385174
rect 311514 349174 312134 384618
rect 311514 348618 311546 349174
rect 312102 348618 312134 349174
rect 311514 313174 312134 348618
rect 311514 312618 311546 313174
rect 312102 312618 312134 313174
rect 311514 277174 312134 312618
rect 311514 276618 311546 277174
rect 312102 276618 312134 277174
rect 311514 241174 312134 276618
rect 311514 240618 311546 241174
rect 312102 240618 312134 241174
rect 311514 205174 312134 240618
rect 311514 204618 311546 205174
rect 312102 204618 312134 205174
rect 311514 169174 312134 204618
rect 311514 168618 311546 169174
rect 312102 168618 312134 169174
rect 311514 133174 312134 168618
rect 311514 132618 311546 133174
rect 312102 132618 312134 133174
rect 311514 97174 312134 132618
rect 311514 96618 311546 97174
rect 312102 96618 312134 97174
rect 311514 61174 312134 96618
rect 311514 60618 311546 61174
rect 312102 60618 312134 61174
rect 311514 25174 312134 60618
rect 311514 24618 311546 25174
rect 312102 24618 312134 25174
rect 311514 -3226 312134 24618
rect 311514 -3782 311546 -3226
rect 312102 -3782 312134 -3226
rect 311514 -3814 312134 -3782
rect 315234 676894 315854 709082
rect 315234 676338 315266 676894
rect 315822 676338 315854 676894
rect 315234 640894 315854 676338
rect 315234 640338 315266 640894
rect 315822 640338 315854 640894
rect 315234 604894 315854 640338
rect 315234 604338 315266 604894
rect 315822 604338 315854 604894
rect 315234 568894 315854 604338
rect 315234 568338 315266 568894
rect 315822 568338 315854 568894
rect 315234 532894 315854 568338
rect 315234 532338 315266 532894
rect 315822 532338 315854 532894
rect 315234 496894 315854 532338
rect 315234 496338 315266 496894
rect 315822 496338 315854 496894
rect 315234 460894 315854 496338
rect 315234 460338 315266 460894
rect 315822 460338 315854 460894
rect 315234 424894 315854 460338
rect 315234 424338 315266 424894
rect 315822 424338 315854 424894
rect 315234 388894 315854 424338
rect 315234 388338 315266 388894
rect 315822 388338 315854 388894
rect 315234 352894 315854 388338
rect 315234 352338 315266 352894
rect 315822 352338 315854 352894
rect 315234 316894 315854 352338
rect 315234 316338 315266 316894
rect 315822 316338 315854 316894
rect 315234 280894 315854 316338
rect 315234 280338 315266 280894
rect 315822 280338 315854 280894
rect 315234 244894 315854 280338
rect 315234 244338 315266 244894
rect 315822 244338 315854 244894
rect 315234 208894 315854 244338
rect 315234 208338 315266 208894
rect 315822 208338 315854 208894
rect 315234 172894 315854 208338
rect 315234 172338 315266 172894
rect 315822 172338 315854 172894
rect 315234 136894 315854 172338
rect 315234 136338 315266 136894
rect 315822 136338 315854 136894
rect 315234 100894 315854 136338
rect 315234 100338 315266 100894
rect 315822 100338 315854 100894
rect 315234 64894 315854 100338
rect 315234 64338 315266 64894
rect 315822 64338 315854 64894
rect 315234 28894 315854 64338
rect 315234 28338 315266 28894
rect 315822 28338 315854 28894
rect 315234 -5146 315854 28338
rect 315234 -5702 315266 -5146
rect 315822 -5702 315854 -5146
rect 315234 -5734 315854 -5702
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710042 336986 710598
rect 337542 710042 337574 710598
rect 333234 708678 333854 709670
rect 333234 708122 333266 708678
rect 333822 708122 333854 708678
rect 329514 706758 330134 707750
rect 329514 706202 329546 706758
rect 330102 706202 330134 706758
rect 318954 680058 318986 680614
rect 319542 680058 319574 680614
rect 318954 644614 319574 680058
rect 318954 644058 318986 644614
rect 319542 644058 319574 644614
rect 318954 608614 319574 644058
rect 318954 608058 318986 608614
rect 319542 608058 319574 608614
rect 318954 572614 319574 608058
rect 318954 572058 318986 572614
rect 319542 572058 319574 572614
rect 318954 536614 319574 572058
rect 318954 536058 318986 536614
rect 319542 536058 319574 536614
rect 318954 500614 319574 536058
rect 318954 500058 318986 500614
rect 319542 500058 319574 500614
rect 318954 464614 319574 500058
rect 318954 464058 318986 464614
rect 319542 464058 319574 464614
rect 318954 428614 319574 464058
rect 318954 428058 318986 428614
rect 319542 428058 319574 428614
rect 318954 392614 319574 428058
rect 318954 392058 318986 392614
rect 319542 392058 319574 392614
rect 318954 356614 319574 392058
rect 318954 356058 318986 356614
rect 319542 356058 319574 356614
rect 318954 320614 319574 356058
rect 318954 320058 318986 320614
rect 319542 320058 319574 320614
rect 318954 284614 319574 320058
rect 318954 284058 318986 284614
rect 319542 284058 319574 284614
rect 318954 248614 319574 284058
rect 318954 248058 318986 248614
rect 319542 248058 319574 248614
rect 318954 212614 319574 248058
rect 318954 212058 318986 212614
rect 319542 212058 319574 212614
rect 318954 176614 319574 212058
rect 318954 176058 318986 176614
rect 319542 176058 319574 176614
rect 318954 140614 319574 176058
rect 318954 140058 318986 140614
rect 319542 140058 319574 140614
rect 318954 104614 319574 140058
rect 318954 104058 318986 104614
rect 319542 104058 319574 104614
rect 318954 68614 319574 104058
rect 318954 68058 318986 68614
rect 319542 68058 319574 68614
rect 318954 32614 319574 68058
rect 318954 32058 318986 32614
rect 319542 32058 319574 32614
rect 300954 -6662 300986 -6106
rect 301542 -6662 301574 -6106
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 704838 326414 705830
rect 325794 704282 325826 704838
rect 326382 704282 326414 704838
rect 325794 687454 326414 704282
rect 325794 686898 325826 687454
rect 326382 686898 326414 687454
rect 325794 651454 326414 686898
rect 325794 650898 325826 651454
rect 326382 650898 326414 651454
rect 325794 615454 326414 650898
rect 325794 614898 325826 615454
rect 326382 614898 326414 615454
rect 325794 579454 326414 614898
rect 325794 578898 325826 579454
rect 326382 578898 326414 579454
rect 325794 543454 326414 578898
rect 325794 542898 325826 543454
rect 326382 542898 326414 543454
rect 325794 507454 326414 542898
rect 325794 506898 325826 507454
rect 326382 506898 326414 507454
rect 325794 471454 326414 506898
rect 325794 470898 325826 471454
rect 326382 470898 326414 471454
rect 325794 435454 326414 470898
rect 325794 434898 325826 435454
rect 326382 434898 326414 435454
rect 325794 399454 326414 434898
rect 325794 398898 325826 399454
rect 326382 398898 326414 399454
rect 325794 363454 326414 398898
rect 325794 362898 325826 363454
rect 326382 362898 326414 363454
rect 325794 327454 326414 362898
rect 325794 326898 325826 327454
rect 326382 326898 326414 327454
rect 325794 291454 326414 326898
rect 325794 290898 325826 291454
rect 326382 290898 326414 291454
rect 325794 255454 326414 290898
rect 325794 254898 325826 255454
rect 326382 254898 326414 255454
rect 325794 219454 326414 254898
rect 325794 218898 325826 219454
rect 326382 218898 326414 219454
rect 325794 183454 326414 218898
rect 325794 182898 325826 183454
rect 326382 182898 326414 183454
rect 325794 147454 326414 182898
rect 325794 146898 325826 147454
rect 326382 146898 326414 147454
rect 325794 111454 326414 146898
rect 325794 110898 325826 111454
rect 326382 110898 326414 111454
rect 325794 75454 326414 110898
rect 325794 74898 325826 75454
rect 326382 74898 326414 75454
rect 325794 39454 326414 74898
rect 325794 38898 325826 39454
rect 326382 38898 326414 39454
rect 325794 3454 326414 38898
rect 325794 2898 325826 3454
rect 326382 2898 326414 3454
rect 325794 -346 326414 2898
rect 325794 -902 325826 -346
rect 326382 -902 326414 -346
rect 325794 -1894 326414 -902
rect 329514 691174 330134 706202
rect 329514 690618 329546 691174
rect 330102 690618 330134 691174
rect 329514 655174 330134 690618
rect 329514 654618 329546 655174
rect 330102 654618 330134 655174
rect 329514 619174 330134 654618
rect 329514 618618 329546 619174
rect 330102 618618 330134 619174
rect 329514 583174 330134 618618
rect 329514 582618 329546 583174
rect 330102 582618 330134 583174
rect 329514 547174 330134 582618
rect 329514 546618 329546 547174
rect 330102 546618 330134 547174
rect 329514 511174 330134 546618
rect 329514 510618 329546 511174
rect 330102 510618 330134 511174
rect 329514 475174 330134 510618
rect 329514 474618 329546 475174
rect 330102 474618 330134 475174
rect 329514 439174 330134 474618
rect 329514 438618 329546 439174
rect 330102 438618 330134 439174
rect 329514 403174 330134 438618
rect 329514 402618 329546 403174
rect 330102 402618 330134 403174
rect 329514 367174 330134 402618
rect 329514 366618 329546 367174
rect 330102 366618 330134 367174
rect 329514 331174 330134 366618
rect 329514 330618 329546 331174
rect 330102 330618 330134 331174
rect 329514 295174 330134 330618
rect 329514 294618 329546 295174
rect 330102 294618 330134 295174
rect 329514 259174 330134 294618
rect 329514 258618 329546 259174
rect 330102 258618 330134 259174
rect 329514 223174 330134 258618
rect 329514 222618 329546 223174
rect 330102 222618 330134 223174
rect 329514 187174 330134 222618
rect 329514 186618 329546 187174
rect 330102 186618 330134 187174
rect 329514 151174 330134 186618
rect 329514 150618 329546 151174
rect 330102 150618 330134 151174
rect 329514 115174 330134 150618
rect 329514 114618 329546 115174
rect 330102 114618 330134 115174
rect 329514 79174 330134 114618
rect 329514 78618 329546 79174
rect 330102 78618 330134 79174
rect 329514 43174 330134 78618
rect 329514 42618 329546 43174
rect 330102 42618 330134 43174
rect 329514 7174 330134 42618
rect 329514 6618 329546 7174
rect 330102 6618 330134 7174
rect 329514 -2266 330134 6618
rect 329514 -2822 329546 -2266
rect 330102 -2822 330134 -2266
rect 329514 -3814 330134 -2822
rect 333234 694894 333854 708122
rect 333234 694338 333266 694894
rect 333822 694338 333854 694894
rect 333234 658894 333854 694338
rect 333234 658338 333266 658894
rect 333822 658338 333854 658894
rect 333234 622894 333854 658338
rect 333234 622338 333266 622894
rect 333822 622338 333854 622894
rect 333234 586894 333854 622338
rect 333234 586338 333266 586894
rect 333822 586338 333854 586894
rect 333234 550894 333854 586338
rect 333234 550338 333266 550894
rect 333822 550338 333854 550894
rect 333234 514894 333854 550338
rect 333234 514338 333266 514894
rect 333822 514338 333854 514894
rect 333234 478894 333854 514338
rect 333234 478338 333266 478894
rect 333822 478338 333854 478894
rect 333234 442894 333854 478338
rect 333234 442338 333266 442894
rect 333822 442338 333854 442894
rect 333234 406894 333854 442338
rect 333234 406338 333266 406894
rect 333822 406338 333854 406894
rect 333234 370894 333854 406338
rect 333234 370338 333266 370894
rect 333822 370338 333854 370894
rect 333234 334894 333854 370338
rect 333234 334338 333266 334894
rect 333822 334338 333854 334894
rect 333234 298894 333854 334338
rect 333234 298338 333266 298894
rect 333822 298338 333854 298894
rect 333234 262894 333854 298338
rect 333234 262338 333266 262894
rect 333822 262338 333854 262894
rect 333234 226894 333854 262338
rect 333234 226338 333266 226894
rect 333822 226338 333854 226894
rect 333234 190894 333854 226338
rect 333234 190338 333266 190894
rect 333822 190338 333854 190894
rect 333234 154894 333854 190338
rect 333234 154338 333266 154894
rect 333822 154338 333854 154894
rect 333234 118894 333854 154338
rect 333234 118338 333266 118894
rect 333822 118338 333854 118894
rect 333234 82894 333854 118338
rect 333234 82338 333266 82894
rect 333822 82338 333854 82894
rect 333234 46894 333854 82338
rect 333234 46338 333266 46894
rect 333822 46338 333854 46894
rect 333234 10894 333854 46338
rect 333234 10338 333266 10894
rect 333822 10338 333854 10894
rect 333234 -4186 333854 10338
rect 333234 -4742 333266 -4186
rect 333822 -4742 333854 -4186
rect 333234 -5734 333854 -4742
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711002 354986 711558
rect 355542 711002 355574 711558
rect 351234 709638 351854 709670
rect 351234 709082 351266 709638
rect 351822 709082 351854 709638
rect 347514 707718 348134 707750
rect 347514 707162 347546 707718
rect 348102 707162 348134 707718
rect 336954 698058 336986 698614
rect 337542 698058 337574 698614
rect 336954 662614 337574 698058
rect 336954 662058 336986 662614
rect 337542 662058 337574 662614
rect 336954 626614 337574 662058
rect 336954 626058 336986 626614
rect 337542 626058 337574 626614
rect 336954 590614 337574 626058
rect 336954 590058 336986 590614
rect 337542 590058 337574 590614
rect 336954 554614 337574 590058
rect 336954 554058 336986 554614
rect 337542 554058 337574 554614
rect 336954 518614 337574 554058
rect 336954 518058 336986 518614
rect 337542 518058 337574 518614
rect 336954 482614 337574 518058
rect 336954 482058 336986 482614
rect 337542 482058 337574 482614
rect 336954 446614 337574 482058
rect 336954 446058 336986 446614
rect 337542 446058 337574 446614
rect 336954 410614 337574 446058
rect 336954 410058 336986 410614
rect 337542 410058 337574 410614
rect 336954 374614 337574 410058
rect 336954 374058 336986 374614
rect 337542 374058 337574 374614
rect 336954 338614 337574 374058
rect 336954 338058 336986 338614
rect 337542 338058 337574 338614
rect 336954 302614 337574 338058
rect 336954 302058 336986 302614
rect 337542 302058 337574 302614
rect 336954 266614 337574 302058
rect 336954 266058 336986 266614
rect 337542 266058 337574 266614
rect 336954 230614 337574 266058
rect 336954 230058 336986 230614
rect 337542 230058 337574 230614
rect 336954 194614 337574 230058
rect 336954 194058 336986 194614
rect 337542 194058 337574 194614
rect 336954 158614 337574 194058
rect 336954 158058 336986 158614
rect 337542 158058 337574 158614
rect 336954 122614 337574 158058
rect 336954 122058 336986 122614
rect 337542 122058 337574 122614
rect 336954 86614 337574 122058
rect 336954 86058 336986 86614
rect 337542 86058 337574 86614
rect 336954 50614 337574 86058
rect 336954 50058 336986 50614
rect 337542 50058 337574 50614
rect 336954 14614 337574 50058
rect 336954 14058 336986 14614
rect 337542 14058 337574 14614
rect 318954 -7622 318986 -7066
rect 319542 -7622 319574 -7066
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 705798 344414 705830
rect 343794 705242 343826 705798
rect 344382 705242 344414 705798
rect 343794 669454 344414 705242
rect 343794 668898 343826 669454
rect 344382 668898 344414 669454
rect 343794 633454 344414 668898
rect 343794 632898 343826 633454
rect 344382 632898 344414 633454
rect 343794 597454 344414 632898
rect 343794 596898 343826 597454
rect 344382 596898 344414 597454
rect 343794 561454 344414 596898
rect 343794 560898 343826 561454
rect 344382 560898 344414 561454
rect 343794 525454 344414 560898
rect 343794 524898 343826 525454
rect 344382 524898 344414 525454
rect 343794 489454 344414 524898
rect 343794 488898 343826 489454
rect 344382 488898 344414 489454
rect 343794 453454 344414 488898
rect 343794 452898 343826 453454
rect 344382 452898 344414 453454
rect 343794 417454 344414 452898
rect 343794 416898 343826 417454
rect 344382 416898 344414 417454
rect 343794 381454 344414 416898
rect 343794 380898 343826 381454
rect 344382 380898 344414 381454
rect 343794 345454 344414 380898
rect 343794 344898 343826 345454
rect 344382 344898 344414 345454
rect 343794 309454 344414 344898
rect 343794 308898 343826 309454
rect 344382 308898 344414 309454
rect 343794 273454 344414 308898
rect 343794 272898 343826 273454
rect 344382 272898 344414 273454
rect 343794 237454 344414 272898
rect 343794 236898 343826 237454
rect 344382 236898 344414 237454
rect 343794 201454 344414 236898
rect 343794 200898 343826 201454
rect 344382 200898 344414 201454
rect 343794 165454 344414 200898
rect 343794 164898 343826 165454
rect 344382 164898 344414 165454
rect 343794 129454 344414 164898
rect 343794 128898 343826 129454
rect 344382 128898 344414 129454
rect 343794 93454 344414 128898
rect 343794 92898 343826 93454
rect 344382 92898 344414 93454
rect 343794 57454 344414 92898
rect 343794 56898 343826 57454
rect 344382 56898 344414 57454
rect 343794 21454 344414 56898
rect 343794 20898 343826 21454
rect 344382 20898 344414 21454
rect 343794 -1306 344414 20898
rect 343794 -1862 343826 -1306
rect 344382 -1862 344414 -1306
rect 343794 -1894 344414 -1862
rect 347514 673174 348134 707162
rect 347514 672618 347546 673174
rect 348102 672618 348134 673174
rect 347514 637174 348134 672618
rect 347514 636618 347546 637174
rect 348102 636618 348134 637174
rect 347514 601174 348134 636618
rect 347514 600618 347546 601174
rect 348102 600618 348134 601174
rect 347514 565174 348134 600618
rect 347514 564618 347546 565174
rect 348102 564618 348134 565174
rect 347514 529174 348134 564618
rect 347514 528618 347546 529174
rect 348102 528618 348134 529174
rect 347514 493174 348134 528618
rect 347514 492618 347546 493174
rect 348102 492618 348134 493174
rect 347514 457174 348134 492618
rect 347514 456618 347546 457174
rect 348102 456618 348134 457174
rect 347514 421174 348134 456618
rect 347514 420618 347546 421174
rect 348102 420618 348134 421174
rect 347514 385174 348134 420618
rect 347514 384618 347546 385174
rect 348102 384618 348134 385174
rect 347514 349174 348134 384618
rect 347514 348618 347546 349174
rect 348102 348618 348134 349174
rect 347514 313174 348134 348618
rect 347514 312618 347546 313174
rect 348102 312618 348134 313174
rect 347514 277174 348134 312618
rect 347514 276618 347546 277174
rect 348102 276618 348134 277174
rect 347514 241174 348134 276618
rect 347514 240618 347546 241174
rect 348102 240618 348134 241174
rect 347514 205174 348134 240618
rect 347514 204618 347546 205174
rect 348102 204618 348134 205174
rect 347514 169174 348134 204618
rect 347514 168618 347546 169174
rect 348102 168618 348134 169174
rect 347514 133174 348134 168618
rect 347514 132618 347546 133174
rect 348102 132618 348134 133174
rect 347514 97174 348134 132618
rect 347514 96618 347546 97174
rect 348102 96618 348134 97174
rect 347514 61174 348134 96618
rect 347514 60618 347546 61174
rect 348102 60618 348134 61174
rect 347514 25174 348134 60618
rect 347514 24618 347546 25174
rect 348102 24618 348134 25174
rect 347514 -3226 348134 24618
rect 347514 -3782 347546 -3226
rect 348102 -3782 348134 -3226
rect 347514 -3814 348134 -3782
rect 351234 676894 351854 709082
rect 351234 676338 351266 676894
rect 351822 676338 351854 676894
rect 351234 640894 351854 676338
rect 351234 640338 351266 640894
rect 351822 640338 351854 640894
rect 351234 604894 351854 640338
rect 351234 604338 351266 604894
rect 351822 604338 351854 604894
rect 351234 568894 351854 604338
rect 351234 568338 351266 568894
rect 351822 568338 351854 568894
rect 351234 532894 351854 568338
rect 351234 532338 351266 532894
rect 351822 532338 351854 532894
rect 351234 496894 351854 532338
rect 351234 496338 351266 496894
rect 351822 496338 351854 496894
rect 351234 460894 351854 496338
rect 351234 460338 351266 460894
rect 351822 460338 351854 460894
rect 351234 424894 351854 460338
rect 351234 424338 351266 424894
rect 351822 424338 351854 424894
rect 351234 388894 351854 424338
rect 351234 388338 351266 388894
rect 351822 388338 351854 388894
rect 351234 352894 351854 388338
rect 351234 352338 351266 352894
rect 351822 352338 351854 352894
rect 351234 316894 351854 352338
rect 351234 316338 351266 316894
rect 351822 316338 351854 316894
rect 351234 280894 351854 316338
rect 351234 280338 351266 280894
rect 351822 280338 351854 280894
rect 351234 244894 351854 280338
rect 351234 244338 351266 244894
rect 351822 244338 351854 244894
rect 351234 208894 351854 244338
rect 351234 208338 351266 208894
rect 351822 208338 351854 208894
rect 351234 172894 351854 208338
rect 351234 172338 351266 172894
rect 351822 172338 351854 172894
rect 351234 136894 351854 172338
rect 351234 136338 351266 136894
rect 351822 136338 351854 136894
rect 351234 100894 351854 136338
rect 351234 100338 351266 100894
rect 351822 100338 351854 100894
rect 351234 64894 351854 100338
rect 351234 64338 351266 64894
rect 351822 64338 351854 64894
rect 351234 28894 351854 64338
rect 351234 28338 351266 28894
rect 351822 28338 351854 28894
rect 351234 -5146 351854 28338
rect 351234 -5702 351266 -5146
rect 351822 -5702 351854 -5146
rect 351234 -5734 351854 -5702
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710042 372986 710598
rect 373542 710042 373574 710598
rect 369234 708678 369854 709670
rect 369234 708122 369266 708678
rect 369822 708122 369854 708678
rect 365514 706758 366134 707750
rect 365514 706202 365546 706758
rect 366102 706202 366134 706758
rect 354954 680058 354986 680614
rect 355542 680058 355574 680614
rect 354954 644614 355574 680058
rect 354954 644058 354986 644614
rect 355542 644058 355574 644614
rect 354954 608614 355574 644058
rect 354954 608058 354986 608614
rect 355542 608058 355574 608614
rect 354954 572614 355574 608058
rect 354954 572058 354986 572614
rect 355542 572058 355574 572614
rect 354954 536614 355574 572058
rect 354954 536058 354986 536614
rect 355542 536058 355574 536614
rect 354954 500614 355574 536058
rect 354954 500058 354986 500614
rect 355542 500058 355574 500614
rect 354954 464614 355574 500058
rect 354954 464058 354986 464614
rect 355542 464058 355574 464614
rect 354954 428614 355574 464058
rect 354954 428058 354986 428614
rect 355542 428058 355574 428614
rect 354954 392614 355574 428058
rect 354954 392058 354986 392614
rect 355542 392058 355574 392614
rect 354954 356614 355574 392058
rect 354954 356058 354986 356614
rect 355542 356058 355574 356614
rect 354954 320614 355574 356058
rect 354954 320058 354986 320614
rect 355542 320058 355574 320614
rect 354954 284614 355574 320058
rect 354954 284058 354986 284614
rect 355542 284058 355574 284614
rect 354954 248614 355574 284058
rect 354954 248058 354986 248614
rect 355542 248058 355574 248614
rect 354954 212614 355574 248058
rect 354954 212058 354986 212614
rect 355542 212058 355574 212614
rect 354954 176614 355574 212058
rect 354954 176058 354986 176614
rect 355542 176058 355574 176614
rect 354954 140614 355574 176058
rect 354954 140058 354986 140614
rect 355542 140058 355574 140614
rect 354954 104614 355574 140058
rect 354954 104058 354986 104614
rect 355542 104058 355574 104614
rect 354954 68614 355574 104058
rect 354954 68058 354986 68614
rect 355542 68058 355574 68614
rect 354954 32614 355574 68058
rect 354954 32058 354986 32614
rect 355542 32058 355574 32614
rect 336954 -6662 336986 -6106
rect 337542 -6662 337574 -6106
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 704838 362414 705830
rect 361794 704282 361826 704838
rect 362382 704282 362414 704838
rect 361794 687454 362414 704282
rect 361794 686898 361826 687454
rect 362382 686898 362414 687454
rect 361794 651454 362414 686898
rect 361794 650898 361826 651454
rect 362382 650898 362414 651454
rect 361794 615454 362414 650898
rect 361794 614898 361826 615454
rect 362382 614898 362414 615454
rect 361794 579454 362414 614898
rect 361794 578898 361826 579454
rect 362382 578898 362414 579454
rect 361794 543454 362414 578898
rect 361794 542898 361826 543454
rect 362382 542898 362414 543454
rect 361794 507454 362414 542898
rect 361794 506898 361826 507454
rect 362382 506898 362414 507454
rect 361794 471454 362414 506898
rect 361794 470898 361826 471454
rect 362382 470898 362414 471454
rect 361794 435454 362414 470898
rect 361794 434898 361826 435454
rect 362382 434898 362414 435454
rect 361794 399454 362414 434898
rect 361794 398898 361826 399454
rect 362382 398898 362414 399454
rect 361794 363454 362414 398898
rect 361794 362898 361826 363454
rect 362382 362898 362414 363454
rect 361794 327454 362414 362898
rect 361794 326898 361826 327454
rect 362382 326898 362414 327454
rect 361794 291454 362414 326898
rect 361794 290898 361826 291454
rect 362382 290898 362414 291454
rect 361794 255454 362414 290898
rect 361794 254898 361826 255454
rect 362382 254898 362414 255454
rect 361794 219454 362414 254898
rect 361794 218898 361826 219454
rect 362382 218898 362414 219454
rect 361794 183454 362414 218898
rect 361794 182898 361826 183454
rect 362382 182898 362414 183454
rect 361794 147454 362414 182898
rect 361794 146898 361826 147454
rect 362382 146898 362414 147454
rect 361794 111454 362414 146898
rect 361794 110898 361826 111454
rect 362382 110898 362414 111454
rect 361794 75454 362414 110898
rect 361794 74898 361826 75454
rect 362382 74898 362414 75454
rect 361794 39454 362414 74898
rect 361794 38898 361826 39454
rect 362382 38898 362414 39454
rect 361794 3454 362414 38898
rect 361794 2898 361826 3454
rect 362382 2898 362414 3454
rect 361794 -346 362414 2898
rect 361794 -902 361826 -346
rect 362382 -902 362414 -346
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690618 365546 691174
rect 366102 690618 366134 691174
rect 365514 655174 366134 690618
rect 365514 654618 365546 655174
rect 366102 654618 366134 655174
rect 365514 619174 366134 654618
rect 365514 618618 365546 619174
rect 366102 618618 366134 619174
rect 365514 583174 366134 618618
rect 365514 582618 365546 583174
rect 366102 582618 366134 583174
rect 365514 547174 366134 582618
rect 365514 546618 365546 547174
rect 366102 546618 366134 547174
rect 365514 511174 366134 546618
rect 365514 510618 365546 511174
rect 366102 510618 366134 511174
rect 365514 475174 366134 510618
rect 365514 474618 365546 475174
rect 366102 474618 366134 475174
rect 365514 439174 366134 474618
rect 365514 438618 365546 439174
rect 366102 438618 366134 439174
rect 365514 403174 366134 438618
rect 365514 402618 365546 403174
rect 366102 402618 366134 403174
rect 365514 367174 366134 402618
rect 365514 366618 365546 367174
rect 366102 366618 366134 367174
rect 365514 331174 366134 366618
rect 365514 330618 365546 331174
rect 366102 330618 366134 331174
rect 365514 295174 366134 330618
rect 365514 294618 365546 295174
rect 366102 294618 366134 295174
rect 365514 259174 366134 294618
rect 365514 258618 365546 259174
rect 366102 258618 366134 259174
rect 365514 223174 366134 258618
rect 365514 222618 365546 223174
rect 366102 222618 366134 223174
rect 365514 187174 366134 222618
rect 365514 186618 365546 187174
rect 366102 186618 366134 187174
rect 365514 151174 366134 186618
rect 365514 150618 365546 151174
rect 366102 150618 366134 151174
rect 365514 115174 366134 150618
rect 365514 114618 365546 115174
rect 366102 114618 366134 115174
rect 365514 79174 366134 114618
rect 365514 78618 365546 79174
rect 366102 78618 366134 79174
rect 365514 43174 366134 78618
rect 365514 42618 365546 43174
rect 366102 42618 366134 43174
rect 365514 7174 366134 42618
rect 365514 6618 365546 7174
rect 366102 6618 366134 7174
rect 365514 -2266 366134 6618
rect 365514 -2822 365546 -2266
rect 366102 -2822 366134 -2266
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694338 369266 694894
rect 369822 694338 369854 694894
rect 369234 658894 369854 694338
rect 369234 658338 369266 658894
rect 369822 658338 369854 658894
rect 369234 622894 369854 658338
rect 369234 622338 369266 622894
rect 369822 622338 369854 622894
rect 369234 586894 369854 622338
rect 369234 586338 369266 586894
rect 369822 586338 369854 586894
rect 369234 550894 369854 586338
rect 369234 550338 369266 550894
rect 369822 550338 369854 550894
rect 369234 514894 369854 550338
rect 369234 514338 369266 514894
rect 369822 514338 369854 514894
rect 369234 478894 369854 514338
rect 369234 478338 369266 478894
rect 369822 478338 369854 478894
rect 369234 442894 369854 478338
rect 369234 442338 369266 442894
rect 369822 442338 369854 442894
rect 369234 406894 369854 442338
rect 369234 406338 369266 406894
rect 369822 406338 369854 406894
rect 369234 370894 369854 406338
rect 369234 370338 369266 370894
rect 369822 370338 369854 370894
rect 369234 334894 369854 370338
rect 369234 334338 369266 334894
rect 369822 334338 369854 334894
rect 369234 298894 369854 334338
rect 369234 298338 369266 298894
rect 369822 298338 369854 298894
rect 369234 262894 369854 298338
rect 369234 262338 369266 262894
rect 369822 262338 369854 262894
rect 369234 226894 369854 262338
rect 369234 226338 369266 226894
rect 369822 226338 369854 226894
rect 369234 190894 369854 226338
rect 369234 190338 369266 190894
rect 369822 190338 369854 190894
rect 369234 154894 369854 190338
rect 369234 154338 369266 154894
rect 369822 154338 369854 154894
rect 369234 118894 369854 154338
rect 369234 118338 369266 118894
rect 369822 118338 369854 118894
rect 369234 82894 369854 118338
rect 369234 82338 369266 82894
rect 369822 82338 369854 82894
rect 369234 46894 369854 82338
rect 369234 46338 369266 46894
rect 369822 46338 369854 46894
rect 369234 10894 369854 46338
rect 369234 10338 369266 10894
rect 369822 10338 369854 10894
rect 369234 -4186 369854 10338
rect 369234 -4742 369266 -4186
rect 369822 -4742 369854 -4186
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711002 390986 711558
rect 391542 711002 391574 711558
rect 387234 709638 387854 709670
rect 387234 709082 387266 709638
rect 387822 709082 387854 709638
rect 383514 707718 384134 707750
rect 383514 707162 383546 707718
rect 384102 707162 384134 707718
rect 372954 698058 372986 698614
rect 373542 698058 373574 698614
rect 372954 662614 373574 698058
rect 372954 662058 372986 662614
rect 373542 662058 373574 662614
rect 372954 626614 373574 662058
rect 372954 626058 372986 626614
rect 373542 626058 373574 626614
rect 372954 590614 373574 626058
rect 372954 590058 372986 590614
rect 373542 590058 373574 590614
rect 372954 554614 373574 590058
rect 372954 554058 372986 554614
rect 373542 554058 373574 554614
rect 372954 518614 373574 554058
rect 372954 518058 372986 518614
rect 373542 518058 373574 518614
rect 372954 482614 373574 518058
rect 372954 482058 372986 482614
rect 373542 482058 373574 482614
rect 372954 446614 373574 482058
rect 372954 446058 372986 446614
rect 373542 446058 373574 446614
rect 372954 410614 373574 446058
rect 372954 410058 372986 410614
rect 373542 410058 373574 410614
rect 372954 374614 373574 410058
rect 372954 374058 372986 374614
rect 373542 374058 373574 374614
rect 372954 338614 373574 374058
rect 372954 338058 372986 338614
rect 373542 338058 373574 338614
rect 372954 302614 373574 338058
rect 372954 302058 372986 302614
rect 373542 302058 373574 302614
rect 372954 266614 373574 302058
rect 372954 266058 372986 266614
rect 373542 266058 373574 266614
rect 372954 230614 373574 266058
rect 372954 230058 372986 230614
rect 373542 230058 373574 230614
rect 372954 194614 373574 230058
rect 372954 194058 372986 194614
rect 373542 194058 373574 194614
rect 372954 158614 373574 194058
rect 372954 158058 372986 158614
rect 373542 158058 373574 158614
rect 372954 122614 373574 158058
rect 372954 122058 372986 122614
rect 373542 122058 373574 122614
rect 372954 86614 373574 122058
rect 372954 86058 372986 86614
rect 373542 86058 373574 86614
rect 372954 50614 373574 86058
rect 372954 50058 372986 50614
rect 373542 50058 373574 50614
rect 372954 14614 373574 50058
rect 372954 14058 372986 14614
rect 373542 14058 373574 14614
rect 354954 -7622 354986 -7066
rect 355542 -7622 355574 -7066
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705242 379826 705798
rect 380382 705242 380414 705798
rect 379794 669454 380414 705242
rect 379794 668898 379826 669454
rect 380382 668898 380414 669454
rect 379794 633454 380414 668898
rect 379794 632898 379826 633454
rect 380382 632898 380414 633454
rect 379794 597454 380414 632898
rect 379794 596898 379826 597454
rect 380382 596898 380414 597454
rect 379794 561454 380414 596898
rect 379794 560898 379826 561454
rect 380382 560898 380414 561454
rect 379794 525454 380414 560898
rect 379794 524898 379826 525454
rect 380382 524898 380414 525454
rect 379794 489454 380414 524898
rect 379794 488898 379826 489454
rect 380382 488898 380414 489454
rect 379794 453454 380414 488898
rect 379794 452898 379826 453454
rect 380382 452898 380414 453454
rect 379794 417454 380414 452898
rect 379794 416898 379826 417454
rect 380382 416898 380414 417454
rect 379794 381454 380414 416898
rect 379794 380898 379826 381454
rect 380382 380898 380414 381454
rect 379794 345454 380414 380898
rect 379794 344898 379826 345454
rect 380382 344898 380414 345454
rect 379794 309454 380414 344898
rect 379794 308898 379826 309454
rect 380382 308898 380414 309454
rect 379794 273454 380414 308898
rect 379794 272898 379826 273454
rect 380382 272898 380414 273454
rect 379794 237454 380414 272898
rect 379794 236898 379826 237454
rect 380382 236898 380414 237454
rect 379794 201454 380414 236898
rect 379794 200898 379826 201454
rect 380382 200898 380414 201454
rect 379794 165454 380414 200898
rect 379794 164898 379826 165454
rect 380382 164898 380414 165454
rect 379794 129454 380414 164898
rect 379794 128898 379826 129454
rect 380382 128898 380414 129454
rect 379794 93454 380414 128898
rect 379794 92898 379826 93454
rect 380382 92898 380414 93454
rect 379794 57454 380414 92898
rect 379794 56898 379826 57454
rect 380382 56898 380414 57454
rect 379794 21454 380414 56898
rect 379794 20898 379826 21454
rect 380382 20898 380414 21454
rect 379794 -1306 380414 20898
rect 379794 -1862 379826 -1306
rect 380382 -1862 380414 -1306
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672618 383546 673174
rect 384102 672618 384134 673174
rect 383514 637174 384134 672618
rect 383514 636618 383546 637174
rect 384102 636618 384134 637174
rect 383514 601174 384134 636618
rect 383514 600618 383546 601174
rect 384102 600618 384134 601174
rect 383514 565174 384134 600618
rect 383514 564618 383546 565174
rect 384102 564618 384134 565174
rect 383514 529174 384134 564618
rect 383514 528618 383546 529174
rect 384102 528618 384134 529174
rect 383514 493174 384134 528618
rect 383514 492618 383546 493174
rect 384102 492618 384134 493174
rect 383514 457174 384134 492618
rect 383514 456618 383546 457174
rect 384102 456618 384134 457174
rect 383514 421174 384134 456618
rect 383514 420618 383546 421174
rect 384102 420618 384134 421174
rect 383514 385174 384134 420618
rect 383514 384618 383546 385174
rect 384102 384618 384134 385174
rect 383514 349174 384134 384618
rect 383514 348618 383546 349174
rect 384102 348618 384134 349174
rect 383514 313174 384134 348618
rect 383514 312618 383546 313174
rect 384102 312618 384134 313174
rect 383514 277174 384134 312618
rect 383514 276618 383546 277174
rect 384102 276618 384134 277174
rect 383514 241174 384134 276618
rect 383514 240618 383546 241174
rect 384102 240618 384134 241174
rect 383514 205174 384134 240618
rect 383514 204618 383546 205174
rect 384102 204618 384134 205174
rect 383514 169174 384134 204618
rect 383514 168618 383546 169174
rect 384102 168618 384134 169174
rect 383514 133174 384134 168618
rect 383514 132618 383546 133174
rect 384102 132618 384134 133174
rect 383514 97174 384134 132618
rect 383514 96618 383546 97174
rect 384102 96618 384134 97174
rect 383514 61174 384134 96618
rect 383514 60618 383546 61174
rect 384102 60618 384134 61174
rect 383514 25174 384134 60618
rect 383514 24618 383546 25174
rect 384102 24618 384134 25174
rect 383514 -3226 384134 24618
rect 383514 -3782 383546 -3226
rect 384102 -3782 384134 -3226
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676338 387266 676894
rect 387822 676338 387854 676894
rect 387234 640894 387854 676338
rect 387234 640338 387266 640894
rect 387822 640338 387854 640894
rect 387234 604894 387854 640338
rect 387234 604338 387266 604894
rect 387822 604338 387854 604894
rect 387234 568894 387854 604338
rect 387234 568338 387266 568894
rect 387822 568338 387854 568894
rect 387234 532894 387854 568338
rect 387234 532338 387266 532894
rect 387822 532338 387854 532894
rect 387234 496894 387854 532338
rect 387234 496338 387266 496894
rect 387822 496338 387854 496894
rect 387234 460894 387854 496338
rect 387234 460338 387266 460894
rect 387822 460338 387854 460894
rect 387234 424894 387854 460338
rect 387234 424338 387266 424894
rect 387822 424338 387854 424894
rect 387234 388894 387854 424338
rect 387234 388338 387266 388894
rect 387822 388338 387854 388894
rect 387234 352894 387854 388338
rect 387234 352338 387266 352894
rect 387822 352338 387854 352894
rect 387234 316894 387854 352338
rect 387234 316338 387266 316894
rect 387822 316338 387854 316894
rect 387234 280894 387854 316338
rect 387234 280338 387266 280894
rect 387822 280338 387854 280894
rect 387234 244894 387854 280338
rect 387234 244338 387266 244894
rect 387822 244338 387854 244894
rect 387234 208894 387854 244338
rect 387234 208338 387266 208894
rect 387822 208338 387854 208894
rect 387234 172894 387854 208338
rect 387234 172338 387266 172894
rect 387822 172338 387854 172894
rect 387234 136894 387854 172338
rect 387234 136338 387266 136894
rect 387822 136338 387854 136894
rect 387234 100894 387854 136338
rect 387234 100338 387266 100894
rect 387822 100338 387854 100894
rect 387234 64894 387854 100338
rect 387234 64338 387266 64894
rect 387822 64338 387854 64894
rect 387234 28894 387854 64338
rect 387234 28338 387266 28894
rect 387822 28338 387854 28894
rect 387234 -5146 387854 28338
rect 387234 -5702 387266 -5146
rect 387822 -5702 387854 -5146
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710042 408986 710598
rect 409542 710042 409574 710598
rect 405234 708678 405854 709670
rect 405234 708122 405266 708678
rect 405822 708122 405854 708678
rect 401514 706758 402134 707750
rect 401514 706202 401546 706758
rect 402102 706202 402134 706758
rect 390954 680058 390986 680614
rect 391542 680058 391574 680614
rect 390954 644614 391574 680058
rect 390954 644058 390986 644614
rect 391542 644058 391574 644614
rect 390954 608614 391574 644058
rect 390954 608058 390986 608614
rect 391542 608058 391574 608614
rect 390954 572614 391574 608058
rect 390954 572058 390986 572614
rect 391542 572058 391574 572614
rect 390954 536614 391574 572058
rect 390954 536058 390986 536614
rect 391542 536058 391574 536614
rect 390954 500614 391574 536058
rect 390954 500058 390986 500614
rect 391542 500058 391574 500614
rect 390954 464614 391574 500058
rect 390954 464058 390986 464614
rect 391542 464058 391574 464614
rect 390954 428614 391574 464058
rect 390954 428058 390986 428614
rect 391542 428058 391574 428614
rect 390954 392614 391574 428058
rect 390954 392058 390986 392614
rect 391542 392058 391574 392614
rect 390954 356614 391574 392058
rect 390954 356058 390986 356614
rect 391542 356058 391574 356614
rect 390954 320614 391574 356058
rect 390954 320058 390986 320614
rect 391542 320058 391574 320614
rect 390954 284614 391574 320058
rect 390954 284058 390986 284614
rect 391542 284058 391574 284614
rect 390954 248614 391574 284058
rect 390954 248058 390986 248614
rect 391542 248058 391574 248614
rect 390954 212614 391574 248058
rect 390954 212058 390986 212614
rect 391542 212058 391574 212614
rect 390954 176614 391574 212058
rect 390954 176058 390986 176614
rect 391542 176058 391574 176614
rect 390954 140614 391574 176058
rect 390954 140058 390986 140614
rect 391542 140058 391574 140614
rect 390954 104614 391574 140058
rect 390954 104058 390986 104614
rect 391542 104058 391574 104614
rect 390954 68614 391574 104058
rect 390954 68058 390986 68614
rect 391542 68058 391574 68614
rect 390954 32614 391574 68058
rect 390954 32058 390986 32614
rect 391542 32058 391574 32614
rect 372954 -6662 372986 -6106
rect 373542 -6662 373574 -6106
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704282 397826 704838
rect 398382 704282 398414 704838
rect 397794 687454 398414 704282
rect 397794 686898 397826 687454
rect 398382 686898 398414 687454
rect 397794 651454 398414 686898
rect 397794 650898 397826 651454
rect 398382 650898 398414 651454
rect 397794 615454 398414 650898
rect 397794 614898 397826 615454
rect 398382 614898 398414 615454
rect 397794 579454 398414 614898
rect 397794 578898 397826 579454
rect 398382 578898 398414 579454
rect 397794 543454 398414 578898
rect 397794 542898 397826 543454
rect 398382 542898 398414 543454
rect 397794 507454 398414 542898
rect 397794 506898 397826 507454
rect 398382 506898 398414 507454
rect 397794 471454 398414 506898
rect 397794 470898 397826 471454
rect 398382 470898 398414 471454
rect 397794 435454 398414 470898
rect 397794 434898 397826 435454
rect 398382 434898 398414 435454
rect 397794 399454 398414 434898
rect 397794 398898 397826 399454
rect 398382 398898 398414 399454
rect 397794 363454 398414 398898
rect 397794 362898 397826 363454
rect 398382 362898 398414 363454
rect 397794 327454 398414 362898
rect 397794 326898 397826 327454
rect 398382 326898 398414 327454
rect 397794 291454 398414 326898
rect 397794 290898 397826 291454
rect 398382 290898 398414 291454
rect 397794 255454 398414 290898
rect 397794 254898 397826 255454
rect 398382 254898 398414 255454
rect 397794 219454 398414 254898
rect 397794 218898 397826 219454
rect 398382 218898 398414 219454
rect 397794 183454 398414 218898
rect 397794 182898 397826 183454
rect 398382 182898 398414 183454
rect 397794 147454 398414 182898
rect 397794 146898 397826 147454
rect 398382 146898 398414 147454
rect 397794 111454 398414 146898
rect 397794 110898 397826 111454
rect 398382 110898 398414 111454
rect 397794 75454 398414 110898
rect 397794 74898 397826 75454
rect 398382 74898 398414 75454
rect 397794 39454 398414 74898
rect 397794 38898 397826 39454
rect 398382 38898 398414 39454
rect 397794 3454 398414 38898
rect 397794 2898 397826 3454
rect 398382 2898 398414 3454
rect 397794 -346 398414 2898
rect 397794 -902 397826 -346
rect 398382 -902 398414 -346
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690618 401546 691174
rect 402102 690618 402134 691174
rect 401514 655174 402134 690618
rect 401514 654618 401546 655174
rect 402102 654618 402134 655174
rect 401514 619174 402134 654618
rect 401514 618618 401546 619174
rect 402102 618618 402134 619174
rect 401514 583174 402134 618618
rect 401514 582618 401546 583174
rect 402102 582618 402134 583174
rect 401514 547174 402134 582618
rect 401514 546618 401546 547174
rect 402102 546618 402134 547174
rect 401514 511174 402134 546618
rect 401514 510618 401546 511174
rect 402102 510618 402134 511174
rect 401514 475174 402134 510618
rect 401514 474618 401546 475174
rect 402102 474618 402134 475174
rect 401514 439174 402134 474618
rect 401514 438618 401546 439174
rect 402102 438618 402134 439174
rect 401514 403174 402134 438618
rect 401514 402618 401546 403174
rect 402102 402618 402134 403174
rect 401514 367174 402134 402618
rect 401514 366618 401546 367174
rect 402102 366618 402134 367174
rect 401514 331174 402134 366618
rect 401514 330618 401546 331174
rect 402102 330618 402134 331174
rect 401514 295174 402134 330618
rect 401514 294618 401546 295174
rect 402102 294618 402134 295174
rect 401514 259174 402134 294618
rect 401514 258618 401546 259174
rect 402102 258618 402134 259174
rect 401514 223174 402134 258618
rect 401514 222618 401546 223174
rect 402102 222618 402134 223174
rect 401514 187174 402134 222618
rect 401514 186618 401546 187174
rect 402102 186618 402134 187174
rect 401514 151174 402134 186618
rect 401514 150618 401546 151174
rect 402102 150618 402134 151174
rect 401514 115174 402134 150618
rect 401514 114618 401546 115174
rect 402102 114618 402134 115174
rect 401514 79174 402134 114618
rect 401514 78618 401546 79174
rect 402102 78618 402134 79174
rect 401514 43174 402134 78618
rect 401514 42618 401546 43174
rect 402102 42618 402134 43174
rect 401514 7174 402134 42618
rect 401514 6618 401546 7174
rect 402102 6618 402134 7174
rect 401514 -2266 402134 6618
rect 401514 -2822 401546 -2266
rect 402102 -2822 402134 -2266
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694338 405266 694894
rect 405822 694338 405854 694894
rect 405234 658894 405854 694338
rect 405234 658338 405266 658894
rect 405822 658338 405854 658894
rect 405234 622894 405854 658338
rect 405234 622338 405266 622894
rect 405822 622338 405854 622894
rect 405234 586894 405854 622338
rect 405234 586338 405266 586894
rect 405822 586338 405854 586894
rect 405234 550894 405854 586338
rect 405234 550338 405266 550894
rect 405822 550338 405854 550894
rect 405234 514894 405854 550338
rect 405234 514338 405266 514894
rect 405822 514338 405854 514894
rect 405234 478894 405854 514338
rect 405234 478338 405266 478894
rect 405822 478338 405854 478894
rect 405234 442894 405854 478338
rect 405234 442338 405266 442894
rect 405822 442338 405854 442894
rect 405234 406894 405854 442338
rect 405234 406338 405266 406894
rect 405822 406338 405854 406894
rect 405234 370894 405854 406338
rect 405234 370338 405266 370894
rect 405822 370338 405854 370894
rect 405234 334894 405854 370338
rect 405234 334338 405266 334894
rect 405822 334338 405854 334894
rect 405234 298894 405854 334338
rect 405234 298338 405266 298894
rect 405822 298338 405854 298894
rect 405234 262894 405854 298338
rect 405234 262338 405266 262894
rect 405822 262338 405854 262894
rect 405234 226894 405854 262338
rect 405234 226338 405266 226894
rect 405822 226338 405854 226894
rect 405234 190894 405854 226338
rect 405234 190338 405266 190894
rect 405822 190338 405854 190894
rect 405234 154894 405854 190338
rect 405234 154338 405266 154894
rect 405822 154338 405854 154894
rect 405234 118894 405854 154338
rect 405234 118338 405266 118894
rect 405822 118338 405854 118894
rect 405234 82894 405854 118338
rect 405234 82338 405266 82894
rect 405822 82338 405854 82894
rect 405234 46894 405854 82338
rect 405234 46338 405266 46894
rect 405822 46338 405854 46894
rect 405234 10894 405854 46338
rect 405234 10338 405266 10894
rect 405822 10338 405854 10894
rect 405234 -4186 405854 10338
rect 405234 -4742 405266 -4186
rect 405822 -4742 405854 -4186
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711002 426986 711558
rect 427542 711002 427574 711558
rect 423234 709638 423854 709670
rect 423234 709082 423266 709638
rect 423822 709082 423854 709638
rect 419514 707718 420134 707750
rect 419514 707162 419546 707718
rect 420102 707162 420134 707718
rect 408954 698058 408986 698614
rect 409542 698058 409574 698614
rect 408954 662614 409574 698058
rect 408954 662058 408986 662614
rect 409542 662058 409574 662614
rect 408954 626614 409574 662058
rect 408954 626058 408986 626614
rect 409542 626058 409574 626614
rect 408954 590614 409574 626058
rect 408954 590058 408986 590614
rect 409542 590058 409574 590614
rect 408954 554614 409574 590058
rect 408954 554058 408986 554614
rect 409542 554058 409574 554614
rect 408954 518614 409574 554058
rect 408954 518058 408986 518614
rect 409542 518058 409574 518614
rect 408954 482614 409574 518058
rect 408954 482058 408986 482614
rect 409542 482058 409574 482614
rect 408954 446614 409574 482058
rect 408954 446058 408986 446614
rect 409542 446058 409574 446614
rect 408954 410614 409574 446058
rect 408954 410058 408986 410614
rect 409542 410058 409574 410614
rect 408954 374614 409574 410058
rect 408954 374058 408986 374614
rect 409542 374058 409574 374614
rect 408954 338614 409574 374058
rect 408954 338058 408986 338614
rect 409542 338058 409574 338614
rect 408954 302614 409574 338058
rect 408954 302058 408986 302614
rect 409542 302058 409574 302614
rect 408954 266614 409574 302058
rect 408954 266058 408986 266614
rect 409542 266058 409574 266614
rect 408954 230614 409574 266058
rect 408954 230058 408986 230614
rect 409542 230058 409574 230614
rect 408954 194614 409574 230058
rect 408954 194058 408986 194614
rect 409542 194058 409574 194614
rect 408954 158614 409574 194058
rect 408954 158058 408986 158614
rect 409542 158058 409574 158614
rect 408954 122614 409574 158058
rect 408954 122058 408986 122614
rect 409542 122058 409574 122614
rect 408954 86614 409574 122058
rect 408954 86058 408986 86614
rect 409542 86058 409574 86614
rect 408954 50614 409574 86058
rect 408954 50058 408986 50614
rect 409542 50058 409574 50614
rect 408954 14614 409574 50058
rect 408954 14058 408986 14614
rect 409542 14058 409574 14614
rect 390954 -7622 390986 -7066
rect 391542 -7622 391574 -7066
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705242 415826 705798
rect 416382 705242 416414 705798
rect 415794 669454 416414 705242
rect 415794 668898 415826 669454
rect 416382 668898 416414 669454
rect 415794 633454 416414 668898
rect 415794 632898 415826 633454
rect 416382 632898 416414 633454
rect 415794 597454 416414 632898
rect 415794 596898 415826 597454
rect 416382 596898 416414 597454
rect 415794 561454 416414 596898
rect 415794 560898 415826 561454
rect 416382 560898 416414 561454
rect 415794 525454 416414 560898
rect 415794 524898 415826 525454
rect 416382 524898 416414 525454
rect 415794 489454 416414 524898
rect 415794 488898 415826 489454
rect 416382 488898 416414 489454
rect 415794 453454 416414 488898
rect 415794 452898 415826 453454
rect 416382 452898 416414 453454
rect 415794 417454 416414 452898
rect 415794 416898 415826 417454
rect 416382 416898 416414 417454
rect 415794 381454 416414 416898
rect 415794 380898 415826 381454
rect 416382 380898 416414 381454
rect 415794 345454 416414 380898
rect 415794 344898 415826 345454
rect 416382 344898 416414 345454
rect 415794 309454 416414 344898
rect 415794 308898 415826 309454
rect 416382 308898 416414 309454
rect 415794 273454 416414 308898
rect 415794 272898 415826 273454
rect 416382 272898 416414 273454
rect 415794 237454 416414 272898
rect 415794 236898 415826 237454
rect 416382 236898 416414 237454
rect 415794 201454 416414 236898
rect 415794 200898 415826 201454
rect 416382 200898 416414 201454
rect 415794 165454 416414 200898
rect 415794 164898 415826 165454
rect 416382 164898 416414 165454
rect 415794 129454 416414 164898
rect 415794 128898 415826 129454
rect 416382 128898 416414 129454
rect 415794 93454 416414 128898
rect 415794 92898 415826 93454
rect 416382 92898 416414 93454
rect 415794 57454 416414 92898
rect 415794 56898 415826 57454
rect 416382 56898 416414 57454
rect 415794 21454 416414 56898
rect 415794 20898 415826 21454
rect 416382 20898 416414 21454
rect 415794 -1306 416414 20898
rect 415794 -1862 415826 -1306
rect 416382 -1862 416414 -1306
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672618 419546 673174
rect 420102 672618 420134 673174
rect 419514 637174 420134 672618
rect 419514 636618 419546 637174
rect 420102 636618 420134 637174
rect 419514 601174 420134 636618
rect 419514 600618 419546 601174
rect 420102 600618 420134 601174
rect 419514 565174 420134 600618
rect 419514 564618 419546 565174
rect 420102 564618 420134 565174
rect 419514 529174 420134 564618
rect 419514 528618 419546 529174
rect 420102 528618 420134 529174
rect 419514 493174 420134 528618
rect 419514 492618 419546 493174
rect 420102 492618 420134 493174
rect 419514 457174 420134 492618
rect 419514 456618 419546 457174
rect 420102 456618 420134 457174
rect 419514 421174 420134 456618
rect 419514 420618 419546 421174
rect 420102 420618 420134 421174
rect 419514 385174 420134 420618
rect 419514 384618 419546 385174
rect 420102 384618 420134 385174
rect 419514 349174 420134 384618
rect 419514 348618 419546 349174
rect 420102 348618 420134 349174
rect 419514 313174 420134 348618
rect 419514 312618 419546 313174
rect 420102 312618 420134 313174
rect 419514 277174 420134 312618
rect 419514 276618 419546 277174
rect 420102 276618 420134 277174
rect 419514 241174 420134 276618
rect 419514 240618 419546 241174
rect 420102 240618 420134 241174
rect 419514 205174 420134 240618
rect 419514 204618 419546 205174
rect 420102 204618 420134 205174
rect 419514 169174 420134 204618
rect 419514 168618 419546 169174
rect 420102 168618 420134 169174
rect 419514 133174 420134 168618
rect 419514 132618 419546 133174
rect 420102 132618 420134 133174
rect 419514 97174 420134 132618
rect 419514 96618 419546 97174
rect 420102 96618 420134 97174
rect 419514 61174 420134 96618
rect 419514 60618 419546 61174
rect 420102 60618 420134 61174
rect 419514 25174 420134 60618
rect 419514 24618 419546 25174
rect 420102 24618 420134 25174
rect 419514 -3226 420134 24618
rect 419514 -3782 419546 -3226
rect 420102 -3782 420134 -3226
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676338 423266 676894
rect 423822 676338 423854 676894
rect 423234 640894 423854 676338
rect 423234 640338 423266 640894
rect 423822 640338 423854 640894
rect 423234 604894 423854 640338
rect 423234 604338 423266 604894
rect 423822 604338 423854 604894
rect 423234 568894 423854 604338
rect 423234 568338 423266 568894
rect 423822 568338 423854 568894
rect 423234 532894 423854 568338
rect 423234 532338 423266 532894
rect 423822 532338 423854 532894
rect 423234 496894 423854 532338
rect 423234 496338 423266 496894
rect 423822 496338 423854 496894
rect 423234 460894 423854 496338
rect 423234 460338 423266 460894
rect 423822 460338 423854 460894
rect 423234 424894 423854 460338
rect 423234 424338 423266 424894
rect 423822 424338 423854 424894
rect 423234 388894 423854 424338
rect 423234 388338 423266 388894
rect 423822 388338 423854 388894
rect 423234 352894 423854 388338
rect 423234 352338 423266 352894
rect 423822 352338 423854 352894
rect 423234 316894 423854 352338
rect 423234 316338 423266 316894
rect 423822 316338 423854 316894
rect 423234 280894 423854 316338
rect 423234 280338 423266 280894
rect 423822 280338 423854 280894
rect 423234 244894 423854 280338
rect 423234 244338 423266 244894
rect 423822 244338 423854 244894
rect 423234 208894 423854 244338
rect 423234 208338 423266 208894
rect 423822 208338 423854 208894
rect 423234 172894 423854 208338
rect 423234 172338 423266 172894
rect 423822 172338 423854 172894
rect 423234 136894 423854 172338
rect 423234 136338 423266 136894
rect 423822 136338 423854 136894
rect 423234 100894 423854 136338
rect 423234 100338 423266 100894
rect 423822 100338 423854 100894
rect 423234 64894 423854 100338
rect 423234 64338 423266 64894
rect 423822 64338 423854 64894
rect 423234 28894 423854 64338
rect 423234 28338 423266 28894
rect 423822 28338 423854 28894
rect 423234 -5146 423854 28338
rect 423234 -5702 423266 -5146
rect 423822 -5702 423854 -5146
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710042 444986 710598
rect 445542 710042 445574 710598
rect 441234 708678 441854 709670
rect 441234 708122 441266 708678
rect 441822 708122 441854 708678
rect 437514 706758 438134 707750
rect 437514 706202 437546 706758
rect 438102 706202 438134 706758
rect 426954 680058 426986 680614
rect 427542 680058 427574 680614
rect 426954 644614 427574 680058
rect 426954 644058 426986 644614
rect 427542 644058 427574 644614
rect 426954 608614 427574 644058
rect 426954 608058 426986 608614
rect 427542 608058 427574 608614
rect 426954 572614 427574 608058
rect 426954 572058 426986 572614
rect 427542 572058 427574 572614
rect 426954 536614 427574 572058
rect 426954 536058 426986 536614
rect 427542 536058 427574 536614
rect 426954 500614 427574 536058
rect 426954 500058 426986 500614
rect 427542 500058 427574 500614
rect 426954 464614 427574 500058
rect 426954 464058 426986 464614
rect 427542 464058 427574 464614
rect 426954 428614 427574 464058
rect 426954 428058 426986 428614
rect 427542 428058 427574 428614
rect 426954 392614 427574 428058
rect 426954 392058 426986 392614
rect 427542 392058 427574 392614
rect 426954 356614 427574 392058
rect 426954 356058 426986 356614
rect 427542 356058 427574 356614
rect 426954 320614 427574 356058
rect 426954 320058 426986 320614
rect 427542 320058 427574 320614
rect 426954 284614 427574 320058
rect 426954 284058 426986 284614
rect 427542 284058 427574 284614
rect 426954 248614 427574 284058
rect 426954 248058 426986 248614
rect 427542 248058 427574 248614
rect 426954 212614 427574 248058
rect 426954 212058 426986 212614
rect 427542 212058 427574 212614
rect 426954 176614 427574 212058
rect 426954 176058 426986 176614
rect 427542 176058 427574 176614
rect 426954 140614 427574 176058
rect 426954 140058 426986 140614
rect 427542 140058 427574 140614
rect 426954 104614 427574 140058
rect 426954 104058 426986 104614
rect 427542 104058 427574 104614
rect 426954 68614 427574 104058
rect 426954 68058 426986 68614
rect 427542 68058 427574 68614
rect 426954 32614 427574 68058
rect 426954 32058 426986 32614
rect 427542 32058 427574 32614
rect 408954 -6662 408986 -6106
rect 409542 -6662 409574 -6106
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704282 433826 704838
rect 434382 704282 434414 704838
rect 433794 687454 434414 704282
rect 433794 686898 433826 687454
rect 434382 686898 434414 687454
rect 433794 651454 434414 686898
rect 433794 650898 433826 651454
rect 434382 650898 434414 651454
rect 433794 615454 434414 650898
rect 433794 614898 433826 615454
rect 434382 614898 434414 615454
rect 433794 579454 434414 614898
rect 433794 578898 433826 579454
rect 434382 578898 434414 579454
rect 433794 543454 434414 578898
rect 433794 542898 433826 543454
rect 434382 542898 434414 543454
rect 433794 507454 434414 542898
rect 433794 506898 433826 507454
rect 434382 506898 434414 507454
rect 433794 471454 434414 506898
rect 433794 470898 433826 471454
rect 434382 470898 434414 471454
rect 433794 435454 434414 470898
rect 433794 434898 433826 435454
rect 434382 434898 434414 435454
rect 433794 399454 434414 434898
rect 433794 398898 433826 399454
rect 434382 398898 434414 399454
rect 433794 363454 434414 398898
rect 433794 362898 433826 363454
rect 434382 362898 434414 363454
rect 433794 327454 434414 362898
rect 433794 326898 433826 327454
rect 434382 326898 434414 327454
rect 433794 291454 434414 326898
rect 433794 290898 433826 291454
rect 434382 290898 434414 291454
rect 433794 255454 434414 290898
rect 433794 254898 433826 255454
rect 434382 254898 434414 255454
rect 433794 219454 434414 254898
rect 433794 218898 433826 219454
rect 434382 218898 434414 219454
rect 433794 183454 434414 218898
rect 433794 182898 433826 183454
rect 434382 182898 434414 183454
rect 433794 147454 434414 182898
rect 433794 146898 433826 147454
rect 434382 146898 434414 147454
rect 433794 111454 434414 146898
rect 433794 110898 433826 111454
rect 434382 110898 434414 111454
rect 433794 75454 434414 110898
rect 433794 74898 433826 75454
rect 434382 74898 434414 75454
rect 433794 39454 434414 74898
rect 433794 38898 433826 39454
rect 434382 38898 434414 39454
rect 433794 3454 434414 38898
rect 433794 2898 433826 3454
rect 434382 2898 434414 3454
rect 433794 -346 434414 2898
rect 433794 -902 433826 -346
rect 434382 -902 434414 -346
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690618 437546 691174
rect 438102 690618 438134 691174
rect 437514 655174 438134 690618
rect 437514 654618 437546 655174
rect 438102 654618 438134 655174
rect 437514 619174 438134 654618
rect 437514 618618 437546 619174
rect 438102 618618 438134 619174
rect 437514 583174 438134 618618
rect 437514 582618 437546 583174
rect 438102 582618 438134 583174
rect 437514 547174 438134 582618
rect 437514 546618 437546 547174
rect 438102 546618 438134 547174
rect 437514 511174 438134 546618
rect 437514 510618 437546 511174
rect 438102 510618 438134 511174
rect 437514 475174 438134 510618
rect 437514 474618 437546 475174
rect 438102 474618 438134 475174
rect 437514 439174 438134 474618
rect 437514 438618 437546 439174
rect 438102 438618 438134 439174
rect 437514 403174 438134 438618
rect 437514 402618 437546 403174
rect 438102 402618 438134 403174
rect 437514 367174 438134 402618
rect 437514 366618 437546 367174
rect 438102 366618 438134 367174
rect 437514 331174 438134 366618
rect 437514 330618 437546 331174
rect 438102 330618 438134 331174
rect 437514 295174 438134 330618
rect 437514 294618 437546 295174
rect 438102 294618 438134 295174
rect 437514 259174 438134 294618
rect 437514 258618 437546 259174
rect 438102 258618 438134 259174
rect 437514 223174 438134 258618
rect 437514 222618 437546 223174
rect 438102 222618 438134 223174
rect 437514 187174 438134 222618
rect 437514 186618 437546 187174
rect 438102 186618 438134 187174
rect 437514 151174 438134 186618
rect 437514 150618 437546 151174
rect 438102 150618 438134 151174
rect 437514 115174 438134 150618
rect 437514 114618 437546 115174
rect 438102 114618 438134 115174
rect 437514 79174 438134 114618
rect 437514 78618 437546 79174
rect 438102 78618 438134 79174
rect 437514 43174 438134 78618
rect 437514 42618 437546 43174
rect 438102 42618 438134 43174
rect 437514 7174 438134 42618
rect 437514 6618 437546 7174
rect 438102 6618 438134 7174
rect 437514 -2266 438134 6618
rect 437514 -2822 437546 -2266
rect 438102 -2822 438134 -2266
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694338 441266 694894
rect 441822 694338 441854 694894
rect 441234 658894 441854 694338
rect 441234 658338 441266 658894
rect 441822 658338 441854 658894
rect 441234 622894 441854 658338
rect 441234 622338 441266 622894
rect 441822 622338 441854 622894
rect 441234 586894 441854 622338
rect 441234 586338 441266 586894
rect 441822 586338 441854 586894
rect 441234 550894 441854 586338
rect 441234 550338 441266 550894
rect 441822 550338 441854 550894
rect 441234 514894 441854 550338
rect 441234 514338 441266 514894
rect 441822 514338 441854 514894
rect 441234 478894 441854 514338
rect 441234 478338 441266 478894
rect 441822 478338 441854 478894
rect 441234 442894 441854 478338
rect 441234 442338 441266 442894
rect 441822 442338 441854 442894
rect 441234 406894 441854 442338
rect 441234 406338 441266 406894
rect 441822 406338 441854 406894
rect 441234 370894 441854 406338
rect 441234 370338 441266 370894
rect 441822 370338 441854 370894
rect 441234 334894 441854 370338
rect 441234 334338 441266 334894
rect 441822 334338 441854 334894
rect 441234 298894 441854 334338
rect 441234 298338 441266 298894
rect 441822 298338 441854 298894
rect 441234 262894 441854 298338
rect 441234 262338 441266 262894
rect 441822 262338 441854 262894
rect 441234 226894 441854 262338
rect 441234 226338 441266 226894
rect 441822 226338 441854 226894
rect 441234 190894 441854 226338
rect 441234 190338 441266 190894
rect 441822 190338 441854 190894
rect 441234 154894 441854 190338
rect 441234 154338 441266 154894
rect 441822 154338 441854 154894
rect 441234 118894 441854 154338
rect 441234 118338 441266 118894
rect 441822 118338 441854 118894
rect 441234 82894 441854 118338
rect 441234 82338 441266 82894
rect 441822 82338 441854 82894
rect 441234 46894 441854 82338
rect 441234 46338 441266 46894
rect 441822 46338 441854 46894
rect 441234 10894 441854 46338
rect 441234 10338 441266 10894
rect 441822 10338 441854 10894
rect 441234 -4186 441854 10338
rect 441234 -4742 441266 -4186
rect 441822 -4742 441854 -4186
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711002 462986 711558
rect 463542 711002 463574 711558
rect 459234 709638 459854 709670
rect 459234 709082 459266 709638
rect 459822 709082 459854 709638
rect 455514 707718 456134 707750
rect 455514 707162 455546 707718
rect 456102 707162 456134 707718
rect 444954 698058 444986 698614
rect 445542 698058 445574 698614
rect 444954 662614 445574 698058
rect 444954 662058 444986 662614
rect 445542 662058 445574 662614
rect 444954 626614 445574 662058
rect 444954 626058 444986 626614
rect 445542 626058 445574 626614
rect 444954 590614 445574 626058
rect 444954 590058 444986 590614
rect 445542 590058 445574 590614
rect 444954 554614 445574 590058
rect 444954 554058 444986 554614
rect 445542 554058 445574 554614
rect 444954 518614 445574 554058
rect 444954 518058 444986 518614
rect 445542 518058 445574 518614
rect 444954 482614 445574 518058
rect 444954 482058 444986 482614
rect 445542 482058 445574 482614
rect 444954 446614 445574 482058
rect 444954 446058 444986 446614
rect 445542 446058 445574 446614
rect 444954 410614 445574 446058
rect 444954 410058 444986 410614
rect 445542 410058 445574 410614
rect 444954 374614 445574 410058
rect 444954 374058 444986 374614
rect 445542 374058 445574 374614
rect 444954 338614 445574 374058
rect 444954 338058 444986 338614
rect 445542 338058 445574 338614
rect 444954 302614 445574 338058
rect 444954 302058 444986 302614
rect 445542 302058 445574 302614
rect 444954 266614 445574 302058
rect 444954 266058 444986 266614
rect 445542 266058 445574 266614
rect 444954 230614 445574 266058
rect 444954 230058 444986 230614
rect 445542 230058 445574 230614
rect 444954 194614 445574 230058
rect 444954 194058 444986 194614
rect 445542 194058 445574 194614
rect 444954 158614 445574 194058
rect 444954 158058 444986 158614
rect 445542 158058 445574 158614
rect 444954 122614 445574 158058
rect 444954 122058 444986 122614
rect 445542 122058 445574 122614
rect 444954 86614 445574 122058
rect 444954 86058 444986 86614
rect 445542 86058 445574 86614
rect 444954 50614 445574 86058
rect 444954 50058 444986 50614
rect 445542 50058 445574 50614
rect 444954 14614 445574 50058
rect 444954 14058 444986 14614
rect 445542 14058 445574 14614
rect 426954 -7622 426986 -7066
rect 427542 -7622 427574 -7066
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705242 451826 705798
rect 452382 705242 452414 705798
rect 451794 669454 452414 705242
rect 451794 668898 451826 669454
rect 452382 668898 452414 669454
rect 451794 633454 452414 668898
rect 451794 632898 451826 633454
rect 452382 632898 452414 633454
rect 451794 597454 452414 632898
rect 451794 596898 451826 597454
rect 452382 596898 452414 597454
rect 451794 561454 452414 596898
rect 451794 560898 451826 561454
rect 452382 560898 452414 561454
rect 451794 525454 452414 560898
rect 451794 524898 451826 525454
rect 452382 524898 452414 525454
rect 451794 489454 452414 524898
rect 451794 488898 451826 489454
rect 452382 488898 452414 489454
rect 451794 453454 452414 488898
rect 451794 452898 451826 453454
rect 452382 452898 452414 453454
rect 451794 417454 452414 452898
rect 451794 416898 451826 417454
rect 452382 416898 452414 417454
rect 451794 381454 452414 416898
rect 451794 380898 451826 381454
rect 452382 380898 452414 381454
rect 451794 345454 452414 380898
rect 451794 344898 451826 345454
rect 452382 344898 452414 345454
rect 451794 309454 452414 344898
rect 451794 308898 451826 309454
rect 452382 308898 452414 309454
rect 451794 273454 452414 308898
rect 451794 272898 451826 273454
rect 452382 272898 452414 273454
rect 451794 237454 452414 272898
rect 451794 236898 451826 237454
rect 452382 236898 452414 237454
rect 451794 201454 452414 236898
rect 451794 200898 451826 201454
rect 452382 200898 452414 201454
rect 451794 165454 452414 200898
rect 451794 164898 451826 165454
rect 452382 164898 452414 165454
rect 451794 129454 452414 164898
rect 451794 128898 451826 129454
rect 452382 128898 452414 129454
rect 451794 93454 452414 128898
rect 451794 92898 451826 93454
rect 452382 92898 452414 93454
rect 451794 57454 452414 92898
rect 451794 56898 451826 57454
rect 452382 56898 452414 57454
rect 451794 21454 452414 56898
rect 451794 20898 451826 21454
rect 452382 20898 452414 21454
rect 451794 -1306 452414 20898
rect 451794 -1862 451826 -1306
rect 452382 -1862 452414 -1306
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672618 455546 673174
rect 456102 672618 456134 673174
rect 455514 637174 456134 672618
rect 455514 636618 455546 637174
rect 456102 636618 456134 637174
rect 455514 601174 456134 636618
rect 455514 600618 455546 601174
rect 456102 600618 456134 601174
rect 455514 565174 456134 600618
rect 455514 564618 455546 565174
rect 456102 564618 456134 565174
rect 455514 529174 456134 564618
rect 455514 528618 455546 529174
rect 456102 528618 456134 529174
rect 455514 493174 456134 528618
rect 455514 492618 455546 493174
rect 456102 492618 456134 493174
rect 455514 457174 456134 492618
rect 455514 456618 455546 457174
rect 456102 456618 456134 457174
rect 455514 421174 456134 456618
rect 455514 420618 455546 421174
rect 456102 420618 456134 421174
rect 455514 385174 456134 420618
rect 455514 384618 455546 385174
rect 456102 384618 456134 385174
rect 455514 349174 456134 384618
rect 455514 348618 455546 349174
rect 456102 348618 456134 349174
rect 455514 313174 456134 348618
rect 455514 312618 455546 313174
rect 456102 312618 456134 313174
rect 455514 277174 456134 312618
rect 455514 276618 455546 277174
rect 456102 276618 456134 277174
rect 455514 241174 456134 276618
rect 455514 240618 455546 241174
rect 456102 240618 456134 241174
rect 455514 205174 456134 240618
rect 455514 204618 455546 205174
rect 456102 204618 456134 205174
rect 455514 169174 456134 204618
rect 455514 168618 455546 169174
rect 456102 168618 456134 169174
rect 455514 133174 456134 168618
rect 455514 132618 455546 133174
rect 456102 132618 456134 133174
rect 455514 97174 456134 132618
rect 455514 96618 455546 97174
rect 456102 96618 456134 97174
rect 455514 61174 456134 96618
rect 455514 60618 455546 61174
rect 456102 60618 456134 61174
rect 455514 25174 456134 60618
rect 455514 24618 455546 25174
rect 456102 24618 456134 25174
rect 455514 -3226 456134 24618
rect 455514 -3782 455546 -3226
rect 456102 -3782 456134 -3226
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676338 459266 676894
rect 459822 676338 459854 676894
rect 459234 640894 459854 676338
rect 459234 640338 459266 640894
rect 459822 640338 459854 640894
rect 459234 604894 459854 640338
rect 459234 604338 459266 604894
rect 459822 604338 459854 604894
rect 459234 568894 459854 604338
rect 459234 568338 459266 568894
rect 459822 568338 459854 568894
rect 459234 532894 459854 568338
rect 459234 532338 459266 532894
rect 459822 532338 459854 532894
rect 459234 496894 459854 532338
rect 459234 496338 459266 496894
rect 459822 496338 459854 496894
rect 459234 460894 459854 496338
rect 459234 460338 459266 460894
rect 459822 460338 459854 460894
rect 459234 424894 459854 460338
rect 459234 424338 459266 424894
rect 459822 424338 459854 424894
rect 459234 388894 459854 424338
rect 459234 388338 459266 388894
rect 459822 388338 459854 388894
rect 459234 352894 459854 388338
rect 459234 352338 459266 352894
rect 459822 352338 459854 352894
rect 459234 316894 459854 352338
rect 459234 316338 459266 316894
rect 459822 316338 459854 316894
rect 459234 280894 459854 316338
rect 459234 280338 459266 280894
rect 459822 280338 459854 280894
rect 459234 244894 459854 280338
rect 459234 244338 459266 244894
rect 459822 244338 459854 244894
rect 459234 208894 459854 244338
rect 459234 208338 459266 208894
rect 459822 208338 459854 208894
rect 459234 172894 459854 208338
rect 459234 172338 459266 172894
rect 459822 172338 459854 172894
rect 459234 136894 459854 172338
rect 459234 136338 459266 136894
rect 459822 136338 459854 136894
rect 459234 100894 459854 136338
rect 459234 100338 459266 100894
rect 459822 100338 459854 100894
rect 459234 64894 459854 100338
rect 459234 64338 459266 64894
rect 459822 64338 459854 64894
rect 459234 28894 459854 64338
rect 459234 28338 459266 28894
rect 459822 28338 459854 28894
rect 459234 -5146 459854 28338
rect 459234 -5702 459266 -5146
rect 459822 -5702 459854 -5146
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710042 480986 710598
rect 481542 710042 481574 710598
rect 477234 708678 477854 709670
rect 477234 708122 477266 708678
rect 477822 708122 477854 708678
rect 473514 706758 474134 707750
rect 473514 706202 473546 706758
rect 474102 706202 474134 706758
rect 462954 680058 462986 680614
rect 463542 680058 463574 680614
rect 462954 644614 463574 680058
rect 462954 644058 462986 644614
rect 463542 644058 463574 644614
rect 462954 608614 463574 644058
rect 462954 608058 462986 608614
rect 463542 608058 463574 608614
rect 462954 572614 463574 608058
rect 462954 572058 462986 572614
rect 463542 572058 463574 572614
rect 462954 536614 463574 572058
rect 462954 536058 462986 536614
rect 463542 536058 463574 536614
rect 462954 500614 463574 536058
rect 462954 500058 462986 500614
rect 463542 500058 463574 500614
rect 462954 464614 463574 500058
rect 462954 464058 462986 464614
rect 463542 464058 463574 464614
rect 462954 428614 463574 464058
rect 462954 428058 462986 428614
rect 463542 428058 463574 428614
rect 462954 392614 463574 428058
rect 462954 392058 462986 392614
rect 463542 392058 463574 392614
rect 462954 356614 463574 392058
rect 462954 356058 462986 356614
rect 463542 356058 463574 356614
rect 462954 320614 463574 356058
rect 462954 320058 462986 320614
rect 463542 320058 463574 320614
rect 462954 284614 463574 320058
rect 462954 284058 462986 284614
rect 463542 284058 463574 284614
rect 462954 248614 463574 284058
rect 462954 248058 462986 248614
rect 463542 248058 463574 248614
rect 462954 212614 463574 248058
rect 462954 212058 462986 212614
rect 463542 212058 463574 212614
rect 462954 176614 463574 212058
rect 462954 176058 462986 176614
rect 463542 176058 463574 176614
rect 462954 140614 463574 176058
rect 462954 140058 462986 140614
rect 463542 140058 463574 140614
rect 462954 104614 463574 140058
rect 462954 104058 462986 104614
rect 463542 104058 463574 104614
rect 462954 68614 463574 104058
rect 462954 68058 462986 68614
rect 463542 68058 463574 68614
rect 462954 32614 463574 68058
rect 462954 32058 462986 32614
rect 463542 32058 463574 32614
rect 444954 -6662 444986 -6106
rect 445542 -6662 445574 -6106
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704282 469826 704838
rect 470382 704282 470414 704838
rect 469794 687454 470414 704282
rect 469794 686898 469826 687454
rect 470382 686898 470414 687454
rect 469794 651454 470414 686898
rect 469794 650898 469826 651454
rect 470382 650898 470414 651454
rect 469794 615454 470414 650898
rect 469794 614898 469826 615454
rect 470382 614898 470414 615454
rect 469794 579454 470414 614898
rect 469794 578898 469826 579454
rect 470382 578898 470414 579454
rect 469794 543454 470414 578898
rect 469794 542898 469826 543454
rect 470382 542898 470414 543454
rect 469794 507454 470414 542898
rect 469794 506898 469826 507454
rect 470382 506898 470414 507454
rect 469794 471454 470414 506898
rect 469794 470898 469826 471454
rect 470382 470898 470414 471454
rect 469794 435454 470414 470898
rect 469794 434898 469826 435454
rect 470382 434898 470414 435454
rect 469794 399454 470414 434898
rect 469794 398898 469826 399454
rect 470382 398898 470414 399454
rect 469794 363454 470414 398898
rect 469794 362898 469826 363454
rect 470382 362898 470414 363454
rect 469794 327454 470414 362898
rect 469794 326898 469826 327454
rect 470382 326898 470414 327454
rect 469794 291454 470414 326898
rect 469794 290898 469826 291454
rect 470382 290898 470414 291454
rect 469794 255454 470414 290898
rect 469794 254898 469826 255454
rect 470382 254898 470414 255454
rect 469794 219454 470414 254898
rect 469794 218898 469826 219454
rect 470382 218898 470414 219454
rect 469794 183454 470414 218898
rect 469794 182898 469826 183454
rect 470382 182898 470414 183454
rect 469794 147454 470414 182898
rect 469794 146898 469826 147454
rect 470382 146898 470414 147454
rect 469794 111454 470414 146898
rect 469794 110898 469826 111454
rect 470382 110898 470414 111454
rect 469794 75454 470414 110898
rect 469794 74898 469826 75454
rect 470382 74898 470414 75454
rect 469794 39454 470414 74898
rect 469794 38898 469826 39454
rect 470382 38898 470414 39454
rect 469794 3454 470414 38898
rect 469794 2898 469826 3454
rect 470382 2898 470414 3454
rect 469794 -346 470414 2898
rect 469794 -902 469826 -346
rect 470382 -902 470414 -346
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690618 473546 691174
rect 474102 690618 474134 691174
rect 473514 655174 474134 690618
rect 473514 654618 473546 655174
rect 474102 654618 474134 655174
rect 473514 619174 474134 654618
rect 473514 618618 473546 619174
rect 474102 618618 474134 619174
rect 473514 583174 474134 618618
rect 473514 582618 473546 583174
rect 474102 582618 474134 583174
rect 473514 547174 474134 582618
rect 473514 546618 473546 547174
rect 474102 546618 474134 547174
rect 473514 511174 474134 546618
rect 473514 510618 473546 511174
rect 474102 510618 474134 511174
rect 473514 475174 474134 510618
rect 473514 474618 473546 475174
rect 474102 474618 474134 475174
rect 473514 439174 474134 474618
rect 473514 438618 473546 439174
rect 474102 438618 474134 439174
rect 473514 403174 474134 438618
rect 473514 402618 473546 403174
rect 474102 402618 474134 403174
rect 473514 367174 474134 402618
rect 473514 366618 473546 367174
rect 474102 366618 474134 367174
rect 473514 331174 474134 366618
rect 473514 330618 473546 331174
rect 474102 330618 474134 331174
rect 473514 295174 474134 330618
rect 473514 294618 473546 295174
rect 474102 294618 474134 295174
rect 473514 259174 474134 294618
rect 473514 258618 473546 259174
rect 474102 258618 474134 259174
rect 473514 223174 474134 258618
rect 473514 222618 473546 223174
rect 474102 222618 474134 223174
rect 473514 187174 474134 222618
rect 473514 186618 473546 187174
rect 474102 186618 474134 187174
rect 473514 151174 474134 186618
rect 473514 150618 473546 151174
rect 474102 150618 474134 151174
rect 473514 115174 474134 150618
rect 473514 114618 473546 115174
rect 474102 114618 474134 115174
rect 473514 79174 474134 114618
rect 473514 78618 473546 79174
rect 474102 78618 474134 79174
rect 473514 43174 474134 78618
rect 473514 42618 473546 43174
rect 474102 42618 474134 43174
rect 473514 7174 474134 42618
rect 473514 6618 473546 7174
rect 474102 6618 474134 7174
rect 473514 -2266 474134 6618
rect 473514 -2822 473546 -2266
rect 474102 -2822 474134 -2266
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694338 477266 694894
rect 477822 694338 477854 694894
rect 477234 658894 477854 694338
rect 477234 658338 477266 658894
rect 477822 658338 477854 658894
rect 477234 622894 477854 658338
rect 477234 622338 477266 622894
rect 477822 622338 477854 622894
rect 477234 586894 477854 622338
rect 477234 586338 477266 586894
rect 477822 586338 477854 586894
rect 477234 550894 477854 586338
rect 477234 550338 477266 550894
rect 477822 550338 477854 550894
rect 477234 514894 477854 550338
rect 477234 514338 477266 514894
rect 477822 514338 477854 514894
rect 477234 478894 477854 514338
rect 477234 478338 477266 478894
rect 477822 478338 477854 478894
rect 477234 442894 477854 478338
rect 477234 442338 477266 442894
rect 477822 442338 477854 442894
rect 477234 406894 477854 442338
rect 477234 406338 477266 406894
rect 477822 406338 477854 406894
rect 477234 370894 477854 406338
rect 477234 370338 477266 370894
rect 477822 370338 477854 370894
rect 477234 334894 477854 370338
rect 477234 334338 477266 334894
rect 477822 334338 477854 334894
rect 477234 298894 477854 334338
rect 477234 298338 477266 298894
rect 477822 298338 477854 298894
rect 477234 262894 477854 298338
rect 477234 262338 477266 262894
rect 477822 262338 477854 262894
rect 477234 226894 477854 262338
rect 477234 226338 477266 226894
rect 477822 226338 477854 226894
rect 477234 190894 477854 226338
rect 477234 190338 477266 190894
rect 477822 190338 477854 190894
rect 477234 154894 477854 190338
rect 477234 154338 477266 154894
rect 477822 154338 477854 154894
rect 477234 118894 477854 154338
rect 477234 118338 477266 118894
rect 477822 118338 477854 118894
rect 477234 82894 477854 118338
rect 477234 82338 477266 82894
rect 477822 82338 477854 82894
rect 477234 46894 477854 82338
rect 477234 46338 477266 46894
rect 477822 46338 477854 46894
rect 477234 10894 477854 46338
rect 477234 10338 477266 10894
rect 477822 10338 477854 10894
rect 477234 -4186 477854 10338
rect 477234 -4742 477266 -4186
rect 477822 -4742 477854 -4186
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711002 498986 711558
rect 499542 711002 499574 711558
rect 495234 709638 495854 709670
rect 495234 709082 495266 709638
rect 495822 709082 495854 709638
rect 491514 707718 492134 707750
rect 491514 707162 491546 707718
rect 492102 707162 492134 707718
rect 480954 698058 480986 698614
rect 481542 698058 481574 698614
rect 480954 662614 481574 698058
rect 480954 662058 480986 662614
rect 481542 662058 481574 662614
rect 480954 626614 481574 662058
rect 480954 626058 480986 626614
rect 481542 626058 481574 626614
rect 480954 590614 481574 626058
rect 480954 590058 480986 590614
rect 481542 590058 481574 590614
rect 480954 554614 481574 590058
rect 480954 554058 480986 554614
rect 481542 554058 481574 554614
rect 480954 518614 481574 554058
rect 480954 518058 480986 518614
rect 481542 518058 481574 518614
rect 480954 482614 481574 518058
rect 480954 482058 480986 482614
rect 481542 482058 481574 482614
rect 480954 446614 481574 482058
rect 480954 446058 480986 446614
rect 481542 446058 481574 446614
rect 480954 410614 481574 446058
rect 480954 410058 480986 410614
rect 481542 410058 481574 410614
rect 480954 374614 481574 410058
rect 480954 374058 480986 374614
rect 481542 374058 481574 374614
rect 480954 338614 481574 374058
rect 480954 338058 480986 338614
rect 481542 338058 481574 338614
rect 480954 302614 481574 338058
rect 480954 302058 480986 302614
rect 481542 302058 481574 302614
rect 480954 266614 481574 302058
rect 480954 266058 480986 266614
rect 481542 266058 481574 266614
rect 480954 230614 481574 266058
rect 480954 230058 480986 230614
rect 481542 230058 481574 230614
rect 480954 194614 481574 230058
rect 480954 194058 480986 194614
rect 481542 194058 481574 194614
rect 480954 158614 481574 194058
rect 480954 158058 480986 158614
rect 481542 158058 481574 158614
rect 480954 122614 481574 158058
rect 480954 122058 480986 122614
rect 481542 122058 481574 122614
rect 480954 86614 481574 122058
rect 480954 86058 480986 86614
rect 481542 86058 481574 86614
rect 480954 50614 481574 86058
rect 480954 50058 480986 50614
rect 481542 50058 481574 50614
rect 480954 14614 481574 50058
rect 480954 14058 480986 14614
rect 481542 14058 481574 14614
rect 462954 -7622 462986 -7066
rect 463542 -7622 463574 -7066
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705242 487826 705798
rect 488382 705242 488414 705798
rect 487794 669454 488414 705242
rect 487794 668898 487826 669454
rect 488382 668898 488414 669454
rect 487794 633454 488414 668898
rect 487794 632898 487826 633454
rect 488382 632898 488414 633454
rect 487794 597454 488414 632898
rect 487794 596898 487826 597454
rect 488382 596898 488414 597454
rect 487794 561454 488414 596898
rect 487794 560898 487826 561454
rect 488382 560898 488414 561454
rect 487794 525454 488414 560898
rect 487794 524898 487826 525454
rect 488382 524898 488414 525454
rect 487794 489454 488414 524898
rect 487794 488898 487826 489454
rect 488382 488898 488414 489454
rect 487794 453454 488414 488898
rect 487794 452898 487826 453454
rect 488382 452898 488414 453454
rect 487794 417454 488414 452898
rect 487794 416898 487826 417454
rect 488382 416898 488414 417454
rect 487794 381454 488414 416898
rect 487794 380898 487826 381454
rect 488382 380898 488414 381454
rect 487794 345454 488414 380898
rect 487794 344898 487826 345454
rect 488382 344898 488414 345454
rect 487794 309454 488414 344898
rect 487794 308898 487826 309454
rect 488382 308898 488414 309454
rect 487794 273454 488414 308898
rect 487794 272898 487826 273454
rect 488382 272898 488414 273454
rect 487794 237454 488414 272898
rect 487794 236898 487826 237454
rect 488382 236898 488414 237454
rect 487794 201454 488414 236898
rect 487794 200898 487826 201454
rect 488382 200898 488414 201454
rect 487794 165454 488414 200898
rect 487794 164898 487826 165454
rect 488382 164898 488414 165454
rect 487794 129454 488414 164898
rect 487794 128898 487826 129454
rect 488382 128898 488414 129454
rect 487794 93454 488414 128898
rect 487794 92898 487826 93454
rect 488382 92898 488414 93454
rect 487794 57454 488414 92898
rect 487794 56898 487826 57454
rect 488382 56898 488414 57454
rect 487794 21454 488414 56898
rect 487794 20898 487826 21454
rect 488382 20898 488414 21454
rect 487794 -1306 488414 20898
rect 487794 -1862 487826 -1306
rect 488382 -1862 488414 -1306
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672618 491546 673174
rect 492102 672618 492134 673174
rect 491514 637174 492134 672618
rect 491514 636618 491546 637174
rect 492102 636618 492134 637174
rect 491514 601174 492134 636618
rect 491514 600618 491546 601174
rect 492102 600618 492134 601174
rect 491514 565174 492134 600618
rect 491514 564618 491546 565174
rect 492102 564618 492134 565174
rect 491514 529174 492134 564618
rect 491514 528618 491546 529174
rect 492102 528618 492134 529174
rect 491514 493174 492134 528618
rect 491514 492618 491546 493174
rect 492102 492618 492134 493174
rect 491514 457174 492134 492618
rect 491514 456618 491546 457174
rect 492102 456618 492134 457174
rect 491514 421174 492134 456618
rect 491514 420618 491546 421174
rect 492102 420618 492134 421174
rect 491514 385174 492134 420618
rect 491514 384618 491546 385174
rect 492102 384618 492134 385174
rect 491514 349174 492134 384618
rect 491514 348618 491546 349174
rect 492102 348618 492134 349174
rect 491514 313174 492134 348618
rect 491514 312618 491546 313174
rect 492102 312618 492134 313174
rect 491514 277174 492134 312618
rect 491514 276618 491546 277174
rect 492102 276618 492134 277174
rect 491514 241174 492134 276618
rect 491514 240618 491546 241174
rect 492102 240618 492134 241174
rect 491514 205174 492134 240618
rect 491514 204618 491546 205174
rect 492102 204618 492134 205174
rect 491514 169174 492134 204618
rect 491514 168618 491546 169174
rect 492102 168618 492134 169174
rect 491514 133174 492134 168618
rect 491514 132618 491546 133174
rect 492102 132618 492134 133174
rect 491514 97174 492134 132618
rect 491514 96618 491546 97174
rect 492102 96618 492134 97174
rect 491514 61174 492134 96618
rect 491514 60618 491546 61174
rect 492102 60618 492134 61174
rect 491514 25174 492134 60618
rect 491514 24618 491546 25174
rect 492102 24618 492134 25174
rect 491514 -3226 492134 24618
rect 491514 -3782 491546 -3226
rect 492102 -3782 492134 -3226
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676338 495266 676894
rect 495822 676338 495854 676894
rect 495234 640894 495854 676338
rect 495234 640338 495266 640894
rect 495822 640338 495854 640894
rect 495234 604894 495854 640338
rect 495234 604338 495266 604894
rect 495822 604338 495854 604894
rect 495234 568894 495854 604338
rect 495234 568338 495266 568894
rect 495822 568338 495854 568894
rect 495234 532894 495854 568338
rect 495234 532338 495266 532894
rect 495822 532338 495854 532894
rect 495234 496894 495854 532338
rect 495234 496338 495266 496894
rect 495822 496338 495854 496894
rect 495234 460894 495854 496338
rect 495234 460338 495266 460894
rect 495822 460338 495854 460894
rect 495234 424894 495854 460338
rect 495234 424338 495266 424894
rect 495822 424338 495854 424894
rect 495234 388894 495854 424338
rect 495234 388338 495266 388894
rect 495822 388338 495854 388894
rect 495234 352894 495854 388338
rect 495234 352338 495266 352894
rect 495822 352338 495854 352894
rect 495234 316894 495854 352338
rect 495234 316338 495266 316894
rect 495822 316338 495854 316894
rect 495234 280894 495854 316338
rect 495234 280338 495266 280894
rect 495822 280338 495854 280894
rect 495234 244894 495854 280338
rect 495234 244338 495266 244894
rect 495822 244338 495854 244894
rect 495234 208894 495854 244338
rect 495234 208338 495266 208894
rect 495822 208338 495854 208894
rect 495234 172894 495854 208338
rect 495234 172338 495266 172894
rect 495822 172338 495854 172894
rect 495234 136894 495854 172338
rect 495234 136338 495266 136894
rect 495822 136338 495854 136894
rect 495234 100894 495854 136338
rect 495234 100338 495266 100894
rect 495822 100338 495854 100894
rect 495234 64894 495854 100338
rect 495234 64338 495266 64894
rect 495822 64338 495854 64894
rect 495234 28894 495854 64338
rect 495234 28338 495266 28894
rect 495822 28338 495854 28894
rect 495234 -5146 495854 28338
rect 495234 -5702 495266 -5146
rect 495822 -5702 495854 -5146
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710042 516986 710598
rect 517542 710042 517574 710598
rect 513234 708678 513854 709670
rect 513234 708122 513266 708678
rect 513822 708122 513854 708678
rect 509514 706758 510134 707750
rect 509514 706202 509546 706758
rect 510102 706202 510134 706758
rect 498954 680058 498986 680614
rect 499542 680058 499574 680614
rect 498954 644614 499574 680058
rect 498954 644058 498986 644614
rect 499542 644058 499574 644614
rect 498954 608614 499574 644058
rect 498954 608058 498986 608614
rect 499542 608058 499574 608614
rect 498954 572614 499574 608058
rect 498954 572058 498986 572614
rect 499542 572058 499574 572614
rect 498954 536614 499574 572058
rect 498954 536058 498986 536614
rect 499542 536058 499574 536614
rect 498954 500614 499574 536058
rect 498954 500058 498986 500614
rect 499542 500058 499574 500614
rect 498954 464614 499574 500058
rect 498954 464058 498986 464614
rect 499542 464058 499574 464614
rect 498954 428614 499574 464058
rect 498954 428058 498986 428614
rect 499542 428058 499574 428614
rect 498954 392614 499574 428058
rect 498954 392058 498986 392614
rect 499542 392058 499574 392614
rect 498954 356614 499574 392058
rect 498954 356058 498986 356614
rect 499542 356058 499574 356614
rect 498954 320614 499574 356058
rect 498954 320058 498986 320614
rect 499542 320058 499574 320614
rect 498954 284614 499574 320058
rect 498954 284058 498986 284614
rect 499542 284058 499574 284614
rect 498954 248614 499574 284058
rect 498954 248058 498986 248614
rect 499542 248058 499574 248614
rect 498954 212614 499574 248058
rect 498954 212058 498986 212614
rect 499542 212058 499574 212614
rect 498954 176614 499574 212058
rect 498954 176058 498986 176614
rect 499542 176058 499574 176614
rect 498954 140614 499574 176058
rect 498954 140058 498986 140614
rect 499542 140058 499574 140614
rect 498954 104614 499574 140058
rect 498954 104058 498986 104614
rect 499542 104058 499574 104614
rect 498954 68614 499574 104058
rect 498954 68058 498986 68614
rect 499542 68058 499574 68614
rect 498954 32614 499574 68058
rect 498954 32058 498986 32614
rect 499542 32058 499574 32614
rect 480954 -6662 480986 -6106
rect 481542 -6662 481574 -6106
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704282 505826 704838
rect 506382 704282 506414 704838
rect 505794 687454 506414 704282
rect 505794 686898 505826 687454
rect 506382 686898 506414 687454
rect 505794 651454 506414 686898
rect 505794 650898 505826 651454
rect 506382 650898 506414 651454
rect 505794 615454 506414 650898
rect 505794 614898 505826 615454
rect 506382 614898 506414 615454
rect 505794 579454 506414 614898
rect 505794 578898 505826 579454
rect 506382 578898 506414 579454
rect 505794 543454 506414 578898
rect 505794 542898 505826 543454
rect 506382 542898 506414 543454
rect 505794 507454 506414 542898
rect 505794 506898 505826 507454
rect 506382 506898 506414 507454
rect 505794 471454 506414 506898
rect 505794 470898 505826 471454
rect 506382 470898 506414 471454
rect 505794 435454 506414 470898
rect 505794 434898 505826 435454
rect 506382 434898 506414 435454
rect 505794 399454 506414 434898
rect 505794 398898 505826 399454
rect 506382 398898 506414 399454
rect 505794 363454 506414 398898
rect 505794 362898 505826 363454
rect 506382 362898 506414 363454
rect 505794 327454 506414 362898
rect 505794 326898 505826 327454
rect 506382 326898 506414 327454
rect 505794 291454 506414 326898
rect 505794 290898 505826 291454
rect 506382 290898 506414 291454
rect 505794 255454 506414 290898
rect 505794 254898 505826 255454
rect 506382 254898 506414 255454
rect 505794 219454 506414 254898
rect 505794 218898 505826 219454
rect 506382 218898 506414 219454
rect 505794 183454 506414 218898
rect 505794 182898 505826 183454
rect 506382 182898 506414 183454
rect 505794 147454 506414 182898
rect 505794 146898 505826 147454
rect 506382 146898 506414 147454
rect 505794 111454 506414 146898
rect 505794 110898 505826 111454
rect 506382 110898 506414 111454
rect 505794 75454 506414 110898
rect 505794 74898 505826 75454
rect 506382 74898 506414 75454
rect 505794 39454 506414 74898
rect 505794 38898 505826 39454
rect 506382 38898 506414 39454
rect 505794 3454 506414 38898
rect 505794 2898 505826 3454
rect 506382 2898 506414 3454
rect 505794 -346 506414 2898
rect 505794 -902 505826 -346
rect 506382 -902 506414 -346
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690618 509546 691174
rect 510102 690618 510134 691174
rect 509514 655174 510134 690618
rect 509514 654618 509546 655174
rect 510102 654618 510134 655174
rect 509514 619174 510134 654618
rect 509514 618618 509546 619174
rect 510102 618618 510134 619174
rect 509514 583174 510134 618618
rect 509514 582618 509546 583174
rect 510102 582618 510134 583174
rect 509514 547174 510134 582618
rect 509514 546618 509546 547174
rect 510102 546618 510134 547174
rect 509514 511174 510134 546618
rect 509514 510618 509546 511174
rect 510102 510618 510134 511174
rect 509514 475174 510134 510618
rect 509514 474618 509546 475174
rect 510102 474618 510134 475174
rect 509514 439174 510134 474618
rect 509514 438618 509546 439174
rect 510102 438618 510134 439174
rect 509514 403174 510134 438618
rect 509514 402618 509546 403174
rect 510102 402618 510134 403174
rect 509514 367174 510134 402618
rect 509514 366618 509546 367174
rect 510102 366618 510134 367174
rect 509514 331174 510134 366618
rect 509514 330618 509546 331174
rect 510102 330618 510134 331174
rect 509514 295174 510134 330618
rect 509514 294618 509546 295174
rect 510102 294618 510134 295174
rect 509514 259174 510134 294618
rect 509514 258618 509546 259174
rect 510102 258618 510134 259174
rect 509514 223174 510134 258618
rect 509514 222618 509546 223174
rect 510102 222618 510134 223174
rect 509514 187174 510134 222618
rect 509514 186618 509546 187174
rect 510102 186618 510134 187174
rect 509514 151174 510134 186618
rect 509514 150618 509546 151174
rect 510102 150618 510134 151174
rect 509514 115174 510134 150618
rect 509514 114618 509546 115174
rect 510102 114618 510134 115174
rect 509514 79174 510134 114618
rect 509514 78618 509546 79174
rect 510102 78618 510134 79174
rect 509514 43174 510134 78618
rect 509514 42618 509546 43174
rect 510102 42618 510134 43174
rect 509514 7174 510134 42618
rect 509514 6618 509546 7174
rect 510102 6618 510134 7174
rect 509514 -2266 510134 6618
rect 509514 -2822 509546 -2266
rect 510102 -2822 510134 -2266
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694338 513266 694894
rect 513822 694338 513854 694894
rect 513234 658894 513854 694338
rect 513234 658338 513266 658894
rect 513822 658338 513854 658894
rect 513234 622894 513854 658338
rect 513234 622338 513266 622894
rect 513822 622338 513854 622894
rect 513234 586894 513854 622338
rect 513234 586338 513266 586894
rect 513822 586338 513854 586894
rect 513234 550894 513854 586338
rect 513234 550338 513266 550894
rect 513822 550338 513854 550894
rect 513234 514894 513854 550338
rect 513234 514338 513266 514894
rect 513822 514338 513854 514894
rect 513234 478894 513854 514338
rect 513234 478338 513266 478894
rect 513822 478338 513854 478894
rect 513234 442894 513854 478338
rect 513234 442338 513266 442894
rect 513822 442338 513854 442894
rect 513234 406894 513854 442338
rect 513234 406338 513266 406894
rect 513822 406338 513854 406894
rect 513234 370894 513854 406338
rect 513234 370338 513266 370894
rect 513822 370338 513854 370894
rect 513234 334894 513854 370338
rect 513234 334338 513266 334894
rect 513822 334338 513854 334894
rect 513234 298894 513854 334338
rect 513234 298338 513266 298894
rect 513822 298338 513854 298894
rect 513234 262894 513854 298338
rect 513234 262338 513266 262894
rect 513822 262338 513854 262894
rect 513234 226894 513854 262338
rect 513234 226338 513266 226894
rect 513822 226338 513854 226894
rect 513234 190894 513854 226338
rect 513234 190338 513266 190894
rect 513822 190338 513854 190894
rect 513234 154894 513854 190338
rect 513234 154338 513266 154894
rect 513822 154338 513854 154894
rect 513234 118894 513854 154338
rect 513234 118338 513266 118894
rect 513822 118338 513854 118894
rect 513234 82894 513854 118338
rect 513234 82338 513266 82894
rect 513822 82338 513854 82894
rect 513234 46894 513854 82338
rect 513234 46338 513266 46894
rect 513822 46338 513854 46894
rect 513234 10894 513854 46338
rect 513234 10338 513266 10894
rect 513822 10338 513854 10894
rect 513234 -4186 513854 10338
rect 513234 -4742 513266 -4186
rect 513822 -4742 513854 -4186
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711002 534986 711558
rect 535542 711002 535574 711558
rect 531234 709638 531854 709670
rect 531234 709082 531266 709638
rect 531822 709082 531854 709638
rect 527514 707718 528134 707750
rect 527514 707162 527546 707718
rect 528102 707162 528134 707718
rect 516954 698058 516986 698614
rect 517542 698058 517574 698614
rect 516954 662614 517574 698058
rect 516954 662058 516986 662614
rect 517542 662058 517574 662614
rect 516954 626614 517574 662058
rect 516954 626058 516986 626614
rect 517542 626058 517574 626614
rect 516954 590614 517574 626058
rect 516954 590058 516986 590614
rect 517542 590058 517574 590614
rect 516954 554614 517574 590058
rect 516954 554058 516986 554614
rect 517542 554058 517574 554614
rect 516954 518614 517574 554058
rect 516954 518058 516986 518614
rect 517542 518058 517574 518614
rect 516954 482614 517574 518058
rect 516954 482058 516986 482614
rect 517542 482058 517574 482614
rect 516954 446614 517574 482058
rect 516954 446058 516986 446614
rect 517542 446058 517574 446614
rect 516954 410614 517574 446058
rect 516954 410058 516986 410614
rect 517542 410058 517574 410614
rect 516954 374614 517574 410058
rect 516954 374058 516986 374614
rect 517542 374058 517574 374614
rect 516954 338614 517574 374058
rect 516954 338058 516986 338614
rect 517542 338058 517574 338614
rect 516954 302614 517574 338058
rect 516954 302058 516986 302614
rect 517542 302058 517574 302614
rect 516954 266614 517574 302058
rect 516954 266058 516986 266614
rect 517542 266058 517574 266614
rect 516954 230614 517574 266058
rect 516954 230058 516986 230614
rect 517542 230058 517574 230614
rect 516954 194614 517574 230058
rect 516954 194058 516986 194614
rect 517542 194058 517574 194614
rect 516954 158614 517574 194058
rect 516954 158058 516986 158614
rect 517542 158058 517574 158614
rect 516954 122614 517574 158058
rect 516954 122058 516986 122614
rect 517542 122058 517574 122614
rect 516954 86614 517574 122058
rect 516954 86058 516986 86614
rect 517542 86058 517574 86614
rect 516954 50614 517574 86058
rect 516954 50058 516986 50614
rect 517542 50058 517574 50614
rect 516954 14614 517574 50058
rect 516954 14058 516986 14614
rect 517542 14058 517574 14614
rect 498954 -7622 498986 -7066
rect 499542 -7622 499574 -7066
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705242 523826 705798
rect 524382 705242 524414 705798
rect 523794 669454 524414 705242
rect 523794 668898 523826 669454
rect 524382 668898 524414 669454
rect 523794 633454 524414 668898
rect 523794 632898 523826 633454
rect 524382 632898 524414 633454
rect 523794 597454 524414 632898
rect 523794 596898 523826 597454
rect 524382 596898 524414 597454
rect 523794 561454 524414 596898
rect 523794 560898 523826 561454
rect 524382 560898 524414 561454
rect 523794 525454 524414 560898
rect 523794 524898 523826 525454
rect 524382 524898 524414 525454
rect 523794 489454 524414 524898
rect 523794 488898 523826 489454
rect 524382 488898 524414 489454
rect 523794 453454 524414 488898
rect 523794 452898 523826 453454
rect 524382 452898 524414 453454
rect 523794 417454 524414 452898
rect 523794 416898 523826 417454
rect 524382 416898 524414 417454
rect 523794 381454 524414 416898
rect 523794 380898 523826 381454
rect 524382 380898 524414 381454
rect 523794 345454 524414 380898
rect 523794 344898 523826 345454
rect 524382 344898 524414 345454
rect 523794 309454 524414 344898
rect 523794 308898 523826 309454
rect 524382 308898 524414 309454
rect 523794 273454 524414 308898
rect 523794 272898 523826 273454
rect 524382 272898 524414 273454
rect 523794 237454 524414 272898
rect 523794 236898 523826 237454
rect 524382 236898 524414 237454
rect 523794 201454 524414 236898
rect 523794 200898 523826 201454
rect 524382 200898 524414 201454
rect 523794 165454 524414 200898
rect 523794 164898 523826 165454
rect 524382 164898 524414 165454
rect 523794 129454 524414 164898
rect 523794 128898 523826 129454
rect 524382 128898 524414 129454
rect 523794 93454 524414 128898
rect 523794 92898 523826 93454
rect 524382 92898 524414 93454
rect 523794 57454 524414 92898
rect 523794 56898 523826 57454
rect 524382 56898 524414 57454
rect 523794 21454 524414 56898
rect 523794 20898 523826 21454
rect 524382 20898 524414 21454
rect 523794 -1306 524414 20898
rect 523794 -1862 523826 -1306
rect 524382 -1862 524414 -1306
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672618 527546 673174
rect 528102 672618 528134 673174
rect 527514 637174 528134 672618
rect 527514 636618 527546 637174
rect 528102 636618 528134 637174
rect 527514 601174 528134 636618
rect 527514 600618 527546 601174
rect 528102 600618 528134 601174
rect 527514 565174 528134 600618
rect 527514 564618 527546 565174
rect 528102 564618 528134 565174
rect 527514 529174 528134 564618
rect 527514 528618 527546 529174
rect 528102 528618 528134 529174
rect 527514 493174 528134 528618
rect 527514 492618 527546 493174
rect 528102 492618 528134 493174
rect 527514 457174 528134 492618
rect 527514 456618 527546 457174
rect 528102 456618 528134 457174
rect 527514 421174 528134 456618
rect 527514 420618 527546 421174
rect 528102 420618 528134 421174
rect 527514 385174 528134 420618
rect 527514 384618 527546 385174
rect 528102 384618 528134 385174
rect 527514 349174 528134 384618
rect 527514 348618 527546 349174
rect 528102 348618 528134 349174
rect 527514 313174 528134 348618
rect 527514 312618 527546 313174
rect 528102 312618 528134 313174
rect 527514 277174 528134 312618
rect 527514 276618 527546 277174
rect 528102 276618 528134 277174
rect 527514 241174 528134 276618
rect 527514 240618 527546 241174
rect 528102 240618 528134 241174
rect 527514 205174 528134 240618
rect 527514 204618 527546 205174
rect 528102 204618 528134 205174
rect 527514 169174 528134 204618
rect 527514 168618 527546 169174
rect 528102 168618 528134 169174
rect 527514 133174 528134 168618
rect 527514 132618 527546 133174
rect 528102 132618 528134 133174
rect 527514 97174 528134 132618
rect 527514 96618 527546 97174
rect 528102 96618 528134 97174
rect 527514 61174 528134 96618
rect 527514 60618 527546 61174
rect 528102 60618 528134 61174
rect 527514 25174 528134 60618
rect 527514 24618 527546 25174
rect 528102 24618 528134 25174
rect 527514 -3226 528134 24618
rect 527514 -3782 527546 -3226
rect 528102 -3782 528134 -3226
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676338 531266 676894
rect 531822 676338 531854 676894
rect 531234 640894 531854 676338
rect 531234 640338 531266 640894
rect 531822 640338 531854 640894
rect 531234 604894 531854 640338
rect 531234 604338 531266 604894
rect 531822 604338 531854 604894
rect 531234 568894 531854 604338
rect 531234 568338 531266 568894
rect 531822 568338 531854 568894
rect 531234 532894 531854 568338
rect 531234 532338 531266 532894
rect 531822 532338 531854 532894
rect 531234 496894 531854 532338
rect 531234 496338 531266 496894
rect 531822 496338 531854 496894
rect 531234 460894 531854 496338
rect 531234 460338 531266 460894
rect 531822 460338 531854 460894
rect 531234 424894 531854 460338
rect 531234 424338 531266 424894
rect 531822 424338 531854 424894
rect 531234 388894 531854 424338
rect 531234 388338 531266 388894
rect 531822 388338 531854 388894
rect 531234 352894 531854 388338
rect 531234 352338 531266 352894
rect 531822 352338 531854 352894
rect 531234 316894 531854 352338
rect 531234 316338 531266 316894
rect 531822 316338 531854 316894
rect 531234 280894 531854 316338
rect 531234 280338 531266 280894
rect 531822 280338 531854 280894
rect 531234 244894 531854 280338
rect 531234 244338 531266 244894
rect 531822 244338 531854 244894
rect 531234 208894 531854 244338
rect 531234 208338 531266 208894
rect 531822 208338 531854 208894
rect 531234 172894 531854 208338
rect 531234 172338 531266 172894
rect 531822 172338 531854 172894
rect 531234 136894 531854 172338
rect 531234 136338 531266 136894
rect 531822 136338 531854 136894
rect 531234 100894 531854 136338
rect 531234 100338 531266 100894
rect 531822 100338 531854 100894
rect 531234 64894 531854 100338
rect 531234 64338 531266 64894
rect 531822 64338 531854 64894
rect 531234 28894 531854 64338
rect 531234 28338 531266 28894
rect 531822 28338 531854 28894
rect 531234 -5146 531854 28338
rect 531234 -5702 531266 -5146
rect 531822 -5702 531854 -5146
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710042 552986 710598
rect 553542 710042 553574 710598
rect 549234 708678 549854 709670
rect 549234 708122 549266 708678
rect 549822 708122 549854 708678
rect 545514 706758 546134 707750
rect 545514 706202 545546 706758
rect 546102 706202 546134 706758
rect 534954 680058 534986 680614
rect 535542 680058 535574 680614
rect 534954 644614 535574 680058
rect 534954 644058 534986 644614
rect 535542 644058 535574 644614
rect 534954 608614 535574 644058
rect 534954 608058 534986 608614
rect 535542 608058 535574 608614
rect 534954 572614 535574 608058
rect 534954 572058 534986 572614
rect 535542 572058 535574 572614
rect 534954 536614 535574 572058
rect 534954 536058 534986 536614
rect 535542 536058 535574 536614
rect 534954 500614 535574 536058
rect 534954 500058 534986 500614
rect 535542 500058 535574 500614
rect 534954 464614 535574 500058
rect 534954 464058 534986 464614
rect 535542 464058 535574 464614
rect 534954 428614 535574 464058
rect 534954 428058 534986 428614
rect 535542 428058 535574 428614
rect 534954 392614 535574 428058
rect 534954 392058 534986 392614
rect 535542 392058 535574 392614
rect 534954 356614 535574 392058
rect 534954 356058 534986 356614
rect 535542 356058 535574 356614
rect 534954 320614 535574 356058
rect 534954 320058 534986 320614
rect 535542 320058 535574 320614
rect 534954 284614 535574 320058
rect 534954 284058 534986 284614
rect 535542 284058 535574 284614
rect 534954 248614 535574 284058
rect 534954 248058 534986 248614
rect 535542 248058 535574 248614
rect 534954 212614 535574 248058
rect 534954 212058 534986 212614
rect 535542 212058 535574 212614
rect 534954 176614 535574 212058
rect 534954 176058 534986 176614
rect 535542 176058 535574 176614
rect 534954 140614 535574 176058
rect 534954 140058 534986 140614
rect 535542 140058 535574 140614
rect 534954 104614 535574 140058
rect 534954 104058 534986 104614
rect 535542 104058 535574 104614
rect 534954 68614 535574 104058
rect 534954 68058 534986 68614
rect 535542 68058 535574 68614
rect 534954 32614 535574 68058
rect 534954 32058 534986 32614
rect 535542 32058 535574 32614
rect 516954 -6662 516986 -6106
rect 517542 -6662 517574 -6106
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704282 541826 704838
rect 542382 704282 542414 704838
rect 541794 687454 542414 704282
rect 541794 686898 541826 687454
rect 542382 686898 542414 687454
rect 541794 651454 542414 686898
rect 541794 650898 541826 651454
rect 542382 650898 542414 651454
rect 541794 615454 542414 650898
rect 541794 614898 541826 615454
rect 542382 614898 542414 615454
rect 541794 579454 542414 614898
rect 541794 578898 541826 579454
rect 542382 578898 542414 579454
rect 541794 543454 542414 578898
rect 541794 542898 541826 543454
rect 542382 542898 542414 543454
rect 541794 507454 542414 542898
rect 541794 506898 541826 507454
rect 542382 506898 542414 507454
rect 541794 471454 542414 506898
rect 541794 470898 541826 471454
rect 542382 470898 542414 471454
rect 541794 435454 542414 470898
rect 541794 434898 541826 435454
rect 542382 434898 542414 435454
rect 541794 399454 542414 434898
rect 541794 398898 541826 399454
rect 542382 398898 542414 399454
rect 541794 363454 542414 398898
rect 541794 362898 541826 363454
rect 542382 362898 542414 363454
rect 541794 327454 542414 362898
rect 541794 326898 541826 327454
rect 542382 326898 542414 327454
rect 541794 291454 542414 326898
rect 541794 290898 541826 291454
rect 542382 290898 542414 291454
rect 541794 255454 542414 290898
rect 541794 254898 541826 255454
rect 542382 254898 542414 255454
rect 541794 219454 542414 254898
rect 541794 218898 541826 219454
rect 542382 218898 542414 219454
rect 541794 183454 542414 218898
rect 541794 182898 541826 183454
rect 542382 182898 542414 183454
rect 541794 147454 542414 182898
rect 541794 146898 541826 147454
rect 542382 146898 542414 147454
rect 541794 111454 542414 146898
rect 541794 110898 541826 111454
rect 542382 110898 542414 111454
rect 541794 75454 542414 110898
rect 541794 74898 541826 75454
rect 542382 74898 542414 75454
rect 541794 39454 542414 74898
rect 541794 38898 541826 39454
rect 542382 38898 542414 39454
rect 541794 3454 542414 38898
rect 541794 2898 541826 3454
rect 542382 2898 542414 3454
rect 541794 -346 542414 2898
rect 541794 -902 541826 -346
rect 542382 -902 542414 -346
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690618 545546 691174
rect 546102 690618 546134 691174
rect 545514 655174 546134 690618
rect 545514 654618 545546 655174
rect 546102 654618 546134 655174
rect 545514 619174 546134 654618
rect 545514 618618 545546 619174
rect 546102 618618 546134 619174
rect 545514 583174 546134 618618
rect 545514 582618 545546 583174
rect 546102 582618 546134 583174
rect 545514 547174 546134 582618
rect 545514 546618 545546 547174
rect 546102 546618 546134 547174
rect 545514 511174 546134 546618
rect 545514 510618 545546 511174
rect 546102 510618 546134 511174
rect 545514 475174 546134 510618
rect 545514 474618 545546 475174
rect 546102 474618 546134 475174
rect 545514 439174 546134 474618
rect 545514 438618 545546 439174
rect 546102 438618 546134 439174
rect 545514 403174 546134 438618
rect 545514 402618 545546 403174
rect 546102 402618 546134 403174
rect 545514 367174 546134 402618
rect 545514 366618 545546 367174
rect 546102 366618 546134 367174
rect 545514 331174 546134 366618
rect 545514 330618 545546 331174
rect 546102 330618 546134 331174
rect 545514 295174 546134 330618
rect 545514 294618 545546 295174
rect 546102 294618 546134 295174
rect 545514 259174 546134 294618
rect 545514 258618 545546 259174
rect 546102 258618 546134 259174
rect 545514 223174 546134 258618
rect 545514 222618 545546 223174
rect 546102 222618 546134 223174
rect 545514 187174 546134 222618
rect 545514 186618 545546 187174
rect 546102 186618 546134 187174
rect 545514 151174 546134 186618
rect 545514 150618 545546 151174
rect 546102 150618 546134 151174
rect 545514 115174 546134 150618
rect 545514 114618 545546 115174
rect 546102 114618 546134 115174
rect 545514 79174 546134 114618
rect 545514 78618 545546 79174
rect 546102 78618 546134 79174
rect 545514 43174 546134 78618
rect 545514 42618 545546 43174
rect 546102 42618 546134 43174
rect 545514 7174 546134 42618
rect 545514 6618 545546 7174
rect 546102 6618 546134 7174
rect 545514 -2266 546134 6618
rect 545514 -2822 545546 -2266
rect 546102 -2822 546134 -2266
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694338 549266 694894
rect 549822 694338 549854 694894
rect 549234 658894 549854 694338
rect 549234 658338 549266 658894
rect 549822 658338 549854 658894
rect 549234 622894 549854 658338
rect 549234 622338 549266 622894
rect 549822 622338 549854 622894
rect 549234 586894 549854 622338
rect 549234 586338 549266 586894
rect 549822 586338 549854 586894
rect 549234 550894 549854 586338
rect 549234 550338 549266 550894
rect 549822 550338 549854 550894
rect 549234 514894 549854 550338
rect 549234 514338 549266 514894
rect 549822 514338 549854 514894
rect 549234 478894 549854 514338
rect 549234 478338 549266 478894
rect 549822 478338 549854 478894
rect 549234 442894 549854 478338
rect 549234 442338 549266 442894
rect 549822 442338 549854 442894
rect 549234 406894 549854 442338
rect 549234 406338 549266 406894
rect 549822 406338 549854 406894
rect 549234 370894 549854 406338
rect 549234 370338 549266 370894
rect 549822 370338 549854 370894
rect 549234 334894 549854 370338
rect 549234 334338 549266 334894
rect 549822 334338 549854 334894
rect 549234 298894 549854 334338
rect 549234 298338 549266 298894
rect 549822 298338 549854 298894
rect 549234 262894 549854 298338
rect 549234 262338 549266 262894
rect 549822 262338 549854 262894
rect 549234 226894 549854 262338
rect 549234 226338 549266 226894
rect 549822 226338 549854 226894
rect 549234 190894 549854 226338
rect 549234 190338 549266 190894
rect 549822 190338 549854 190894
rect 549234 154894 549854 190338
rect 549234 154338 549266 154894
rect 549822 154338 549854 154894
rect 549234 118894 549854 154338
rect 549234 118338 549266 118894
rect 549822 118338 549854 118894
rect 549234 82894 549854 118338
rect 549234 82338 549266 82894
rect 549822 82338 549854 82894
rect 549234 46894 549854 82338
rect 549234 46338 549266 46894
rect 549822 46338 549854 46894
rect 549234 10894 549854 46338
rect 549234 10338 549266 10894
rect 549822 10338 549854 10894
rect 549234 -4186 549854 10338
rect 549234 -4742 549266 -4186
rect 549822 -4742 549854 -4186
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711002 570986 711558
rect 571542 711002 571574 711558
rect 567234 709638 567854 709670
rect 567234 709082 567266 709638
rect 567822 709082 567854 709638
rect 563514 707718 564134 707750
rect 563514 707162 563546 707718
rect 564102 707162 564134 707718
rect 552954 698058 552986 698614
rect 553542 698058 553574 698614
rect 552954 662614 553574 698058
rect 552954 662058 552986 662614
rect 553542 662058 553574 662614
rect 552954 626614 553574 662058
rect 552954 626058 552986 626614
rect 553542 626058 553574 626614
rect 552954 590614 553574 626058
rect 552954 590058 552986 590614
rect 553542 590058 553574 590614
rect 552954 554614 553574 590058
rect 552954 554058 552986 554614
rect 553542 554058 553574 554614
rect 552954 518614 553574 554058
rect 552954 518058 552986 518614
rect 553542 518058 553574 518614
rect 552954 482614 553574 518058
rect 552954 482058 552986 482614
rect 553542 482058 553574 482614
rect 552954 446614 553574 482058
rect 552954 446058 552986 446614
rect 553542 446058 553574 446614
rect 552954 410614 553574 446058
rect 552954 410058 552986 410614
rect 553542 410058 553574 410614
rect 552954 374614 553574 410058
rect 552954 374058 552986 374614
rect 553542 374058 553574 374614
rect 552954 338614 553574 374058
rect 552954 338058 552986 338614
rect 553542 338058 553574 338614
rect 552954 302614 553574 338058
rect 552954 302058 552986 302614
rect 553542 302058 553574 302614
rect 552954 266614 553574 302058
rect 552954 266058 552986 266614
rect 553542 266058 553574 266614
rect 552954 230614 553574 266058
rect 552954 230058 552986 230614
rect 553542 230058 553574 230614
rect 552954 194614 553574 230058
rect 552954 194058 552986 194614
rect 553542 194058 553574 194614
rect 552954 158614 553574 194058
rect 552954 158058 552986 158614
rect 553542 158058 553574 158614
rect 552954 122614 553574 158058
rect 552954 122058 552986 122614
rect 553542 122058 553574 122614
rect 552954 86614 553574 122058
rect 552954 86058 552986 86614
rect 553542 86058 553574 86614
rect 552954 50614 553574 86058
rect 552954 50058 552986 50614
rect 553542 50058 553574 50614
rect 552954 14614 553574 50058
rect 552954 14058 552986 14614
rect 553542 14058 553574 14614
rect 534954 -7622 534986 -7066
rect 535542 -7622 535574 -7066
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705242 559826 705798
rect 560382 705242 560414 705798
rect 559794 669454 560414 705242
rect 559794 668898 559826 669454
rect 560382 668898 560414 669454
rect 559794 633454 560414 668898
rect 559794 632898 559826 633454
rect 560382 632898 560414 633454
rect 559794 597454 560414 632898
rect 559794 596898 559826 597454
rect 560382 596898 560414 597454
rect 559794 561454 560414 596898
rect 559794 560898 559826 561454
rect 560382 560898 560414 561454
rect 559794 525454 560414 560898
rect 559794 524898 559826 525454
rect 560382 524898 560414 525454
rect 559794 489454 560414 524898
rect 559794 488898 559826 489454
rect 560382 488898 560414 489454
rect 559794 453454 560414 488898
rect 559794 452898 559826 453454
rect 560382 452898 560414 453454
rect 559794 417454 560414 452898
rect 559794 416898 559826 417454
rect 560382 416898 560414 417454
rect 559794 381454 560414 416898
rect 559794 380898 559826 381454
rect 560382 380898 560414 381454
rect 559794 345454 560414 380898
rect 559794 344898 559826 345454
rect 560382 344898 560414 345454
rect 559794 309454 560414 344898
rect 559794 308898 559826 309454
rect 560382 308898 560414 309454
rect 559794 273454 560414 308898
rect 559794 272898 559826 273454
rect 560382 272898 560414 273454
rect 559794 237454 560414 272898
rect 559794 236898 559826 237454
rect 560382 236898 560414 237454
rect 559794 201454 560414 236898
rect 559794 200898 559826 201454
rect 560382 200898 560414 201454
rect 559794 165454 560414 200898
rect 559794 164898 559826 165454
rect 560382 164898 560414 165454
rect 559794 129454 560414 164898
rect 559794 128898 559826 129454
rect 560382 128898 560414 129454
rect 559794 93454 560414 128898
rect 559794 92898 559826 93454
rect 560382 92898 560414 93454
rect 559794 57454 560414 92898
rect 559794 56898 559826 57454
rect 560382 56898 560414 57454
rect 559794 21454 560414 56898
rect 559794 20898 559826 21454
rect 560382 20898 560414 21454
rect 559794 -1306 560414 20898
rect 559794 -1862 559826 -1306
rect 560382 -1862 560414 -1306
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672618 563546 673174
rect 564102 672618 564134 673174
rect 563514 637174 564134 672618
rect 563514 636618 563546 637174
rect 564102 636618 564134 637174
rect 563514 601174 564134 636618
rect 563514 600618 563546 601174
rect 564102 600618 564134 601174
rect 563514 565174 564134 600618
rect 563514 564618 563546 565174
rect 564102 564618 564134 565174
rect 563514 529174 564134 564618
rect 563514 528618 563546 529174
rect 564102 528618 564134 529174
rect 563514 493174 564134 528618
rect 563514 492618 563546 493174
rect 564102 492618 564134 493174
rect 563514 457174 564134 492618
rect 563514 456618 563546 457174
rect 564102 456618 564134 457174
rect 563514 421174 564134 456618
rect 563514 420618 563546 421174
rect 564102 420618 564134 421174
rect 563514 385174 564134 420618
rect 563514 384618 563546 385174
rect 564102 384618 564134 385174
rect 563514 349174 564134 384618
rect 563514 348618 563546 349174
rect 564102 348618 564134 349174
rect 563514 313174 564134 348618
rect 563514 312618 563546 313174
rect 564102 312618 564134 313174
rect 563514 277174 564134 312618
rect 563514 276618 563546 277174
rect 564102 276618 564134 277174
rect 563514 241174 564134 276618
rect 563514 240618 563546 241174
rect 564102 240618 564134 241174
rect 563514 205174 564134 240618
rect 563514 204618 563546 205174
rect 564102 204618 564134 205174
rect 563514 169174 564134 204618
rect 563514 168618 563546 169174
rect 564102 168618 564134 169174
rect 563514 133174 564134 168618
rect 563514 132618 563546 133174
rect 564102 132618 564134 133174
rect 563514 97174 564134 132618
rect 563514 96618 563546 97174
rect 564102 96618 564134 97174
rect 563514 61174 564134 96618
rect 563514 60618 563546 61174
rect 564102 60618 564134 61174
rect 563514 25174 564134 60618
rect 563514 24618 563546 25174
rect 564102 24618 564134 25174
rect 563514 -3226 564134 24618
rect 563514 -3782 563546 -3226
rect 564102 -3782 564134 -3226
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676338 567266 676894
rect 567822 676338 567854 676894
rect 567234 640894 567854 676338
rect 567234 640338 567266 640894
rect 567822 640338 567854 640894
rect 567234 604894 567854 640338
rect 567234 604338 567266 604894
rect 567822 604338 567854 604894
rect 567234 568894 567854 604338
rect 567234 568338 567266 568894
rect 567822 568338 567854 568894
rect 567234 532894 567854 568338
rect 567234 532338 567266 532894
rect 567822 532338 567854 532894
rect 567234 496894 567854 532338
rect 567234 496338 567266 496894
rect 567822 496338 567854 496894
rect 567234 460894 567854 496338
rect 567234 460338 567266 460894
rect 567822 460338 567854 460894
rect 567234 424894 567854 460338
rect 567234 424338 567266 424894
rect 567822 424338 567854 424894
rect 567234 388894 567854 424338
rect 567234 388338 567266 388894
rect 567822 388338 567854 388894
rect 567234 352894 567854 388338
rect 567234 352338 567266 352894
rect 567822 352338 567854 352894
rect 567234 316894 567854 352338
rect 567234 316338 567266 316894
rect 567822 316338 567854 316894
rect 567234 280894 567854 316338
rect 567234 280338 567266 280894
rect 567822 280338 567854 280894
rect 567234 244894 567854 280338
rect 567234 244338 567266 244894
rect 567822 244338 567854 244894
rect 567234 208894 567854 244338
rect 567234 208338 567266 208894
rect 567822 208338 567854 208894
rect 567234 172894 567854 208338
rect 567234 172338 567266 172894
rect 567822 172338 567854 172894
rect 567234 136894 567854 172338
rect 567234 136338 567266 136894
rect 567822 136338 567854 136894
rect 567234 100894 567854 136338
rect 567234 100338 567266 100894
rect 567822 100338 567854 100894
rect 567234 64894 567854 100338
rect 567234 64338 567266 64894
rect 567822 64338 567854 64894
rect 567234 28894 567854 64338
rect 567234 28338 567266 28894
rect 567822 28338 567854 28894
rect 567234 -5146 567854 28338
rect 567234 -5702 567266 -5146
rect 567822 -5702 567854 -5146
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711002 592062 711558
rect 592618 711002 592650 711558
rect 591070 710598 591690 710630
rect 591070 710042 591102 710598
rect 591658 710042 591690 710598
rect 590110 709638 590730 709670
rect 590110 709082 590142 709638
rect 590698 709082 590730 709638
rect 589150 708678 589770 708710
rect 589150 708122 589182 708678
rect 589738 708122 589770 708678
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707162 588222 707718
rect 588778 707162 588810 707718
rect 581514 706202 581546 706758
rect 582102 706202 582134 706758
rect 570954 680058 570986 680614
rect 571542 680058 571574 680614
rect 570954 644614 571574 680058
rect 570954 644058 570986 644614
rect 571542 644058 571574 644614
rect 570954 608614 571574 644058
rect 570954 608058 570986 608614
rect 571542 608058 571574 608614
rect 570954 572614 571574 608058
rect 570954 572058 570986 572614
rect 571542 572058 571574 572614
rect 570954 536614 571574 572058
rect 570954 536058 570986 536614
rect 571542 536058 571574 536614
rect 570954 500614 571574 536058
rect 570954 500058 570986 500614
rect 571542 500058 571574 500614
rect 570954 464614 571574 500058
rect 570954 464058 570986 464614
rect 571542 464058 571574 464614
rect 570954 428614 571574 464058
rect 570954 428058 570986 428614
rect 571542 428058 571574 428614
rect 570954 392614 571574 428058
rect 570954 392058 570986 392614
rect 571542 392058 571574 392614
rect 570954 356614 571574 392058
rect 570954 356058 570986 356614
rect 571542 356058 571574 356614
rect 570954 320614 571574 356058
rect 570954 320058 570986 320614
rect 571542 320058 571574 320614
rect 570954 284614 571574 320058
rect 570954 284058 570986 284614
rect 571542 284058 571574 284614
rect 570954 248614 571574 284058
rect 570954 248058 570986 248614
rect 571542 248058 571574 248614
rect 570954 212614 571574 248058
rect 570954 212058 570986 212614
rect 571542 212058 571574 212614
rect 570954 176614 571574 212058
rect 570954 176058 570986 176614
rect 571542 176058 571574 176614
rect 570954 140614 571574 176058
rect 570954 140058 570986 140614
rect 571542 140058 571574 140614
rect 570954 104614 571574 140058
rect 570954 104058 570986 104614
rect 571542 104058 571574 104614
rect 570954 68614 571574 104058
rect 570954 68058 570986 68614
rect 571542 68058 571574 68614
rect 570954 32614 571574 68058
rect 570954 32058 570986 32614
rect 571542 32058 571574 32614
rect 552954 -6662 552986 -6106
rect 553542 -6662 553574 -6106
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704282 577826 704838
rect 578382 704282 578414 704838
rect 577794 687454 578414 704282
rect 577794 686898 577826 687454
rect 578382 686898 578414 687454
rect 577794 651454 578414 686898
rect 577794 650898 577826 651454
rect 578382 650898 578414 651454
rect 577794 615454 578414 650898
rect 577794 614898 577826 615454
rect 578382 614898 578414 615454
rect 577794 579454 578414 614898
rect 577794 578898 577826 579454
rect 578382 578898 578414 579454
rect 577794 543454 578414 578898
rect 577794 542898 577826 543454
rect 578382 542898 578414 543454
rect 577794 507454 578414 542898
rect 577794 506898 577826 507454
rect 578382 506898 578414 507454
rect 577794 471454 578414 506898
rect 577794 470898 577826 471454
rect 578382 470898 578414 471454
rect 577794 435454 578414 470898
rect 577794 434898 577826 435454
rect 578382 434898 578414 435454
rect 577794 399454 578414 434898
rect 577794 398898 577826 399454
rect 578382 398898 578414 399454
rect 577794 363454 578414 398898
rect 577794 362898 577826 363454
rect 578382 362898 578414 363454
rect 577794 327454 578414 362898
rect 577794 326898 577826 327454
rect 578382 326898 578414 327454
rect 577794 291454 578414 326898
rect 577794 290898 577826 291454
rect 578382 290898 578414 291454
rect 577794 255454 578414 290898
rect 577794 254898 577826 255454
rect 578382 254898 578414 255454
rect 577794 219454 578414 254898
rect 577794 218898 577826 219454
rect 578382 218898 578414 219454
rect 577794 183454 578414 218898
rect 577794 182898 577826 183454
rect 578382 182898 578414 183454
rect 577794 147454 578414 182898
rect 577794 146898 577826 147454
rect 578382 146898 578414 147454
rect 577794 111454 578414 146898
rect 577794 110898 577826 111454
rect 578382 110898 578414 111454
rect 577794 75454 578414 110898
rect 577794 74898 577826 75454
rect 578382 74898 578414 75454
rect 577794 39454 578414 74898
rect 577794 38898 577826 39454
rect 578382 38898 578414 39454
rect 577794 3454 578414 38898
rect 577794 2898 577826 3454
rect 578382 2898 578414 3454
rect 577794 -346 578414 2898
rect 577794 -902 577826 -346
rect 578382 -902 578414 -346
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706202 587262 706758
rect 587818 706202 587850 706758
rect 586270 705798 586890 705830
rect 586270 705242 586302 705798
rect 586858 705242 586890 705798
rect 581514 690618 581546 691174
rect 582102 690618 582134 691174
rect 581514 655174 582134 690618
rect 581514 654618 581546 655174
rect 582102 654618 582134 655174
rect 581514 619174 582134 654618
rect 581514 618618 581546 619174
rect 582102 618618 582134 619174
rect 581514 583174 582134 618618
rect 581514 582618 581546 583174
rect 582102 582618 582134 583174
rect 581514 547174 582134 582618
rect 581514 546618 581546 547174
rect 582102 546618 582134 547174
rect 581514 511174 582134 546618
rect 581514 510618 581546 511174
rect 582102 510618 582134 511174
rect 581514 475174 582134 510618
rect 581514 474618 581546 475174
rect 582102 474618 582134 475174
rect 581514 439174 582134 474618
rect 581514 438618 581546 439174
rect 582102 438618 582134 439174
rect 581514 403174 582134 438618
rect 581514 402618 581546 403174
rect 582102 402618 582134 403174
rect 581514 367174 582134 402618
rect 581514 366618 581546 367174
rect 582102 366618 582134 367174
rect 581514 331174 582134 366618
rect 581514 330618 581546 331174
rect 582102 330618 582134 331174
rect 581514 295174 582134 330618
rect 581514 294618 581546 295174
rect 582102 294618 582134 295174
rect 581514 259174 582134 294618
rect 581514 258618 581546 259174
rect 582102 258618 582134 259174
rect 581514 223174 582134 258618
rect 581514 222618 581546 223174
rect 582102 222618 582134 223174
rect 581514 187174 582134 222618
rect 581514 186618 581546 187174
rect 582102 186618 582134 187174
rect 581514 151174 582134 186618
rect 581514 150618 581546 151174
rect 582102 150618 582134 151174
rect 581514 115174 582134 150618
rect 581514 114618 581546 115174
rect 582102 114618 582134 115174
rect 581514 79174 582134 114618
rect 581514 78618 581546 79174
rect 582102 78618 582134 79174
rect 581514 43174 582134 78618
rect 581514 42618 581546 43174
rect 582102 42618 582134 43174
rect 581514 7174 582134 42618
rect 581514 6618 581546 7174
rect 582102 6618 582134 7174
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704282 585342 704838
rect 585898 704282 585930 704838
rect 585310 687454 585930 704282
rect 585310 686898 585342 687454
rect 585898 686898 585930 687454
rect 585310 651454 585930 686898
rect 585310 650898 585342 651454
rect 585898 650898 585930 651454
rect 585310 615454 585930 650898
rect 585310 614898 585342 615454
rect 585898 614898 585930 615454
rect 585310 579454 585930 614898
rect 585310 578898 585342 579454
rect 585898 578898 585930 579454
rect 585310 543454 585930 578898
rect 585310 542898 585342 543454
rect 585898 542898 585930 543454
rect 585310 507454 585930 542898
rect 585310 506898 585342 507454
rect 585898 506898 585930 507454
rect 585310 471454 585930 506898
rect 585310 470898 585342 471454
rect 585898 470898 585930 471454
rect 585310 435454 585930 470898
rect 585310 434898 585342 435454
rect 585898 434898 585930 435454
rect 585310 399454 585930 434898
rect 585310 398898 585342 399454
rect 585898 398898 585930 399454
rect 585310 363454 585930 398898
rect 585310 362898 585342 363454
rect 585898 362898 585930 363454
rect 585310 327454 585930 362898
rect 585310 326898 585342 327454
rect 585898 326898 585930 327454
rect 585310 291454 585930 326898
rect 585310 290898 585342 291454
rect 585898 290898 585930 291454
rect 585310 255454 585930 290898
rect 585310 254898 585342 255454
rect 585898 254898 585930 255454
rect 585310 219454 585930 254898
rect 585310 218898 585342 219454
rect 585898 218898 585930 219454
rect 585310 183454 585930 218898
rect 585310 182898 585342 183454
rect 585898 182898 585930 183454
rect 585310 147454 585930 182898
rect 585310 146898 585342 147454
rect 585898 146898 585930 147454
rect 585310 111454 585930 146898
rect 585310 110898 585342 111454
rect 585898 110898 585930 111454
rect 585310 75454 585930 110898
rect 585310 74898 585342 75454
rect 585898 74898 585930 75454
rect 585310 39454 585930 74898
rect 585310 38898 585342 39454
rect 585898 38898 585930 39454
rect 585310 3454 585930 38898
rect 585310 2898 585342 3454
rect 585898 2898 585930 3454
rect 585310 -346 585930 2898
rect 585310 -902 585342 -346
rect 585898 -902 585930 -346
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 668898 586302 669454
rect 586858 668898 586890 669454
rect 586270 633454 586890 668898
rect 586270 632898 586302 633454
rect 586858 632898 586890 633454
rect 586270 597454 586890 632898
rect 586270 596898 586302 597454
rect 586858 596898 586890 597454
rect 586270 561454 586890 596898
rect 586270 560898 586302 561454
rect 586858 560898 586890 561454
rect 586270 525454 586890 560898
rect 586270 524898 586302 525454
rect 586858 524898 586890 525454
rect 586270 489454 586890 524898
rect 586270 488898 586302 489454
rect 586858 488898 586890 489454
rect 586270 453454 586890 488898
rect 586270 452898 586302 453454
rect 586858 452898 586890 453454
rect 586270 417454 586890 452898
rect 586270 416898 586302 417454
rect 586858 416898 586890 417454
rect 586270 381454 586890 416898
rect 586270 380898 586302 381454
rect 586858 380898 586890 381454
rect 586270 345454 586890 380898
rect 586270 344898 586302 345454
rect 586858 344898 586890 345454
rect 586270 309454 586890 344898
rect 586270 308898 586302 309454
rect 586858 308898 586890 309454
rect 586270 273454 586890 308898
rect 586270 272898 586302 273454
rect 586858 272898 586890 273454
rect 586270 237454 586890 272898
rect 586270 236898 586302 237454
rect 586858 236898 586890 237454
rect 586270 201454 586890 236898
rect 586270 200898 586302 201454
rect 586858 200898 586890 201454
rect 586270 165454 586890 200898
rect 586270 164898 586302 165454
rect 586858 164898 586890 165454
rect 586270 129454 586890 164898
rect 586270 128898 586302 129454
rect 586858 128898 586890 129454
rect 586270 93454 586890 128898
rect 586270 92898 586302 93454
rect 586858 92898 586890 93454
rect 586270 57454 586890 92898
rect 586270 56898 586302 57454
rect 586858 56898 586890 57454
rect 586270 21454 586890 56898
rect 586270 20898 586302 21454
rect 586858 20898 586890 21454
rect 586270 -1306 586890 20898
rect 586270 -1862 586302 -1306
rect 586858 -1862 586890 -1306
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690618 587262 691174
rect 587818 690618 587850 691174
rect 587230 655174 587850 690618
rect 587230 654618 587262 655174
rect 587818 654618 587850 655174
rect 587230 619174 587850 654618
rect 587230 618618 587262 619174
rect 587818 618618 587850 619174
rect 587230 583174 587850 618618
rect 587230 582618 587262 583174
rect 587818 582618 587850 583174
rect 587230 547174 587850 582618
rect 587230 546618 587262 547174
rect 587818 546618 587850 547174
rect 587230 511174 587850 546618
rect 587230 510618 587262 511174
rect 587818 510618 587850 511174
rect 587230 475174 587850 510618
rect 587230 474618 587262 475174
rect 587818 474618 587850 475174
rect 587230 439174 587850 474618
rect 587230 438618 587262 439174
rect 587818 438618 587850 439174
rect 587230 403174 587850 438618
rect 587230 402618 587262 403174
rect 587818 402618 587850 403174
rect 587230 367174 587850 402618
rect 587230 366618 587262 367174
rect 587818 366618 587850 367174
rect 587230 331174 587850 366618
rect 587230 330618 587262 331174
rect 587818 330618 587850 331174
rect 587230 295174 587850 330618
rect 587230 294618 587262 295174
rect 587818 294618 587850 295174
rect 587230 259174 587850 294618
rect 587230 258618 587262 259174
rect 587818 258618 587850 259174
rect 587230 223174 587850 258618
rect 587230 222618 587262 223174
rect 587818 222618 587850 223174
rect 587230 187174 587850 222618
rect 587230 186618 587262 187174
rect 587818 186618 587850 187174
rect 587230 151174 587850 186618
rect 587230 150618 587262 151174
rect 587818 150618 587850 151174
rect 587230 115174 587850 150618
rect 587230 114618 587262 115174
rect 587818 114618 587850 115174
rect 587230 79174 587850 114618
rect 587230 78618 587262 79174
rect 587818 78618 587850 79174
rect 587230 43174 587850 78618
rect 587230 42618 587262 43174
rect 587818 42618 587850 43174
rect 587230 7174 587850 42618
rect 587230 6618 587262 7174
rect 587818 6618 587850 7174
rect 581514 -2822 581546 -2266
rect 582102 -2822 582134 -2266
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2822 587262 -2266
rect 587818 -2822 587850 -2266
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672618 588222 673174
rect 588778 672618 588810 673174
rect 588190 637174 588810 672618
rect 588190 636618 588222 637174
rect 588778 636618 588810 637174
rect 588190 601174 588810 636618
rect 588190 600618 588222 601174
rect 588778 600618 588810 601174
rect 588190 565174 588810 600618
rect 588190 564618 588222 565174
rect 588778 564618 588810 565174
rect 588190 529174 588810 564618
rect 588190 528618 588222 529174
rect 588778 528618 588810 529174
rect 588190 493174 588810 528618
rect 588190 492618 588222 493174
rect 588778 492618 588810 493174
rect 588190 457174 588810 492618
rect 588190 456618 588222 457174
rect 588778 456618 588810 457174
rect 588190 421174 588810 456618
rect 588190 420618 588222 421174
rect 588778 420618 588810 421174
rect 588190 385174 588810 420618
rect 588190 384618 588222 385174
rect 588778 384618 588810 385174
rect 588190 349174 588810 384618
rect 588190 348618 588222 349174
rect 588778 348618 588810 349174
rect 588190 313174 588810 348618
rect 588190 312618 588222 313174
rect 588778 312618 588810 313174
rect 588190 277174 588810 312618
rect 588190 276618 588222 277174
rect 588778 276618 588810 277174
rect 588190 241174 588810 276618
rect 588190 240618 588222 241174
rect 588778 240618 588810 241174
rect 588190 205174 588810 240618
rect 588190 204618 588222 205174
rect 588778 204618 588810 205174
rect 588190 169174 588810 204618
rect 588190 168618 588222 169174
rect 588778 168618 588810 169174
rect 588190 133174 588810 168618
rect 588190 132618 588222 133174
rect 588778 132618 588810 133174
rect 588190 97174 588810 132618
rect 588190 96618 588222 97174
rect 588778 96618 588810 97174
rect 588190 61174 588810 96618
rect 588190 60618 588222 61174
rect 588778 60618 588810 61174
rect 588190 25174 588810 60618
rect 588190 24618 588222 25174
rect 588778 24618 588810 25174
rect 588190 -3226 588810 24618
rect 588190 -3782 588222 -3226
rect 588778 -3782 588810 -3226
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694338 589182 694894
rect 589738 694338 589770 694894
rect 589150 658894 589770 694338
rect 589150 658338 589182 658894
rect 589738 658338 589770 658894
rect 589150 622894 589770 658338
rect 589150 622338 589182 622894
rect 589738 622338 589770 622894
rect 589150 586894 589770 622338
rect 589150 586338 589182 586894
rect 589738 586338 589770 586894
rect 589150 550894 589770 586338
rect 589150 550338 589182 550894
rect 589738 550338 589770 550894
rect 589150 514894 589770 550338
rect 589150 514338 589182 514894
rect 589738 514338 589770 514894
rect 589150 478894 589770 514338
rect 589150 478338 589182 478894
rect 589738 478338 589770 478894
rect 589150 442894 589770 478338
rect 589150 442338 589182 442894
rect 589738 442338 589770 442894
rect 589150 406894 589770 442338
rect 589150 406338 589182 406894
rect 589738 406338 589770 406894
rect 589150 370894 589770 406338
rect 589150 370338 589182 370894
rect 589738 370338 589770 370894
rect 589150 334894 589770 370338
rect 589150 334338 589182 334894
rect 589738 334338 589770 334894
rect 589150 298894 589770 334338
rect 589150 298338 589182 298894
rect 589738 298338 589770 298894
rect 589150 262894 589770 298338
rect 589150 262338 589182 262894
rect 589738 262338 589770 262894
rect 589150 226894 589770 262338
rect 589150 226338 589182 226894
rect 589738 226338 589770 226894
rect 589150 190894 589770 226338
rect 589150 190338 589182 190894
rect 589738 190338 589770 190894
rect 589150 154894 589770 190338
rect 589150 154338 589182 154894
rect 589738 154338 589770 154894
rect 589150 118894 589770 154338
rect 589150 118338 589182 118894
rect 589738 118338 589770 118894
rect 589150 82894 589770 118338
rect 589150 82338 589182 82894
rect 589738 82338 589770 82894
rect 589150 46894 589770 82338
rect 589150 46338 589182 46894
rect 589738 46338 589770 46894
rect 589150 10894 589770 46338
rect 589150 10338 589182 10894
rect 589738 10338 589770 10894
rect 589150 -4186 589770 10338
rect 589150 -4742 589182 -4186
rect 589738 -4742 589770 -4186
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676338 590142 676894
rect 590698 676338 590730 676894
rect 590110 640894 590730 676338
rect 590110 640338 590142 640894
rect 590698 640338 590730 640894
rect 590110 604894 590730 640338
rect 590110 604338 590142 604894
rect 590698 604338 590730 604894
rect 590110 568894 590730 604338
rect 590110 568338 590142 568894
rect 590698 568338 590730 568894
rect 590110 532894 590730 568338
rect 590110 532338 590142 532894
rect 590698 532338 590730 532894
rect 590110 496894 590730 532338
rect 590110 496338 590142 496894
rect 590698 496338 590730 496894
rect 590110 460894 590730 496338
rect 590110 460338 590142 460894
rect 590698 460338 590730 460894
rect 590110 424894 590730 460338
rect 590110 424338 590142 424894
rect 590698 424338 590730 424894
rect 590110 388894 590730 424338
rect 590110 388338 590142 388894
rect 590698 388338 590730 388894
rect 590110 352894 590730 388338
rect 590110 352338 590142 352894
rect 590698 352338 590730 352894
rect 590110 316894 590730 352338
rect 590110 316338 590142 316894
rect 590698 316338 590730 316894
rect 590110 280894 590730 316338
rect 590110 280338 590142 280894
rect 590698 280338 590730 280894
rect 590110 244894 590730 280338
rect 590110 244338 590142 244894
rect 590698 244338 590730 244894
rect 590110 208894 590730 244338
rect 590110 208338 590142 208894
rect 590698 208338 590730 208894
rect 590110 172894 590730 208338
rect 590110 172338 590142 172894
rect 590698 172338 590730 172894
rect 590110 136894 590730 172338
rect 590110 136338 590142 136894
rect 590698 136338 590730 136894
rect 590110 100894 590730 136338
rect 590110 100338 590142 100894
rect 590698 100338 590730 100894
rect 590110 64894 590730 100338
rect 590110 64338 590142 64894
rect 590698 64338 590730 64894
rect 590110 28894 590730 64338
rect 590110 28338 590142 28894
rect 590698 28338 590730 28894
rect 590110 -5146 590730 28338
rect 590110 -5702 590142 -5146
rect 590698 -5702 590730 -5146
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698058 591102 698614
rect 591658 698058 591690 698614
rect 591070 662614 591690 698058
rect 591070 662058 591102 662614
rect 591658 662058 591690 662614
rect 591070 626614 591690 662058
rect 591070 626058 591102 626614
rect 591658 626058 591690 626614
rect 591070 590614 591690 626058
rect 591070 590058 591102 590614
rect 591658 590058 591690 590614
rect 591070 554614 591690 590058
rect 591070 554058 591102 554614
rect 591658 554058 591690 554614
rect 591070 518614 591690 554058
rect 591070 518058 591102 518614
rect 591658 518058 591690 518614
rect 591070 482614 591690 518058
rect 591070 482058 591102 482614
rect 591658 482058 591690 482614
rect 591070 446614 591690 482058
rect 591070 446058 591102 446614
rect 591658 446058 591690 446614
rect 591070 410614 591690 446058
rect 591070 410058 591102 410614
rect 591658 410058 591690 410614
rect 591070 374614 591690 410058
rect 591070 374058 591102 374614
rect 591658 374058 591690 374614
rect 591070 338614 591690 374058
rect 591070 338058 591102 338614
rect 591658 338058 591690 338614
rect 591070 302614 591690 338058
rect 591070 302058 591102 302614
rect 591658 302058 591690 302614
rect 591070 266614 591690 302058
rect 591070 266058 591102 266614
rect 591658 266058 591690 266614
rect 591070 230614 591690 266058
rect 591070 230058 591102 230614
rect 591658 230058 591690 230614
rect 591070 194614 591690 230058
rect 591070 194058 591102 194614
rect 591658 194058 591690 194614
rect 591070 158614 591690 194058
rect 591070 158058 591102 158614
rect 591658 158058 591690 158614
rect 591070 122614 591690 158058
rect 591070 122058 591102 122614
rect 591658 122058 591690 122614
rect 591070 86614 591690 122058
rect 591070 86058 591102 86614
rect 591658 86058 591690 86614
rect 591070 50614 591690 86058
rect 591070 50058 591102 50614
rect 591658 50058 591690 50614
rect 591070 14614 591690 50058
rect 591070 14058 591102 14614
rect 591658 14058 591690 14614
rect 591070 -6106 591690 14058
rect 591070 -6662 591102 -6106
rect 591658 -6662 591690 -6106
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680058 592062 680614
rect 592618 680058 592650 680614
rect 592030 644614 592650 680058
rect 592030 644058 592062 644614
rect 592618 644058 592650 644614
rect 592030 608614 592650 644058
rect 592030 608058 592062 608614
rect 592618 608058 592650 608614
rect 592030 572614 592650 608058
rect 592030 572058 592062 572614
rect 592618 572058 592650 572614
rect 592030 536614 592650 572058
rect 592030 536058 592062 536614
rect 592618 536058 592650 536614
rect 592030 500614 592650 536058
rect 592030 500058 592062 500614
rect 592618 500058 592650 500614
rect 592030 464614 592650 500058
rect 592030 464058 592062 464614
rect 592618 464058 592650 464614
rect 592030 428614 592650 464058
rect 592030 428058 592062 428614
rect 592618 428058 592650 428614
rect 592030 392614 592650 428058
rect 592030 392058 592062 392614
rect 592618 392058 592650 392614
rect 592030 356614 592650 392058
rect 592030 356058 592062 356614
rect 592618 356058 592650 356614
rect 592030 320614 592650 356058
rect 592030 320058 592062 320614
rect 592618 320058 592650 320614
rect 592030 284614 592650 320058
rect 592030 284058 592062 284614
rect 592618 284058 592650 284614
rect 592030 248614 592650 284058
rect 592030 248058 592062 248614
rect 592618 248058 592650 248614
rect 592030 212614 592650 248058
rect 592030 212058 592062 212614
rect 592618 212058 592650 212614
rect 592030 176614 592650 212058
rect 592030 176058 592062 176614
rect 592618 176058 592650 176614
rect 592030 140614 592650 176058
rect 592030 140058 592062 140614
rect 592618 140058 592650 140614
rect 592030 104614 592650 140058
rect 592030 104058 592062 104614
rect 592618 104058 592650 104614
rect 592030 68614 592650 104058
rect 592030 68058 592062 68614
rect 592618 68058 592650 68614
rect 592030 32614 592650 68058
rect 592030 32058 592062 32614
rect 592618 32058 592650 32614
rect 570954 -7622 570986 -7066
rect 571542 -7622 571574 -7066
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7622 592062 -7066
rect 592618 -7622 592650 -7066
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711002 -8138 711558
rect -8694 680058 -8138 680614
rect -8694 644058 -8138 644614
rect -8694 608058 -8138 608614
rect -8694 572058 -8138 572614
rect -8694 536058 -8138 536614
rect -8694 500058 -8138 500614
rect -8694 464058 -8138 464614
rect -8694 428058 -8138 428614
rect -8694 392058 -8138 392614
rect -8694 356058 -8138 356614
rect -8694 320058 -8138 320614
rect -8694 284058 -8138 284614
rect -8694 248058 -8138 248614
rect -8694 212058 -8138 212614
rect -8694 176058 -8138 176614
rect -8694 140058 -8138 140614
rect -8694 104058 -8138 104614
rect -8694 68058 -8138 68614
rect -8694 32058 -8138 32614
rect -7734 710042 -7178 710598
rect 12986 710042 13542 710598
rect -7734 698058 -7178 698614
rect -7734 662058 -7178 662614
rect -7734 626058 -7178 626614
rect -7734 590058 -7178 590614
rect -7734 554058 -7178 554614
rect -7734 518058 -7178 518614
rect -7734 482058 -7178 482614
rect -7734 446058 -7178 446614
rect -7734 410058 -7178 410614
rect -7734 374058 -7178 374614
rect -7734 338058 -7178 338614
rect -7734 302058 -7178 302614
rect -7734 266058 -7178 266614
rect -7734 230058 -7178 230614
rect -7734 194058 -7178 194614
rect -7734 158058 -7178 158614
rect -7734 122058 -7178 122614
rect -7734 86058 -7178 86614
rect -7734 50058 -7178 50614
rect -7734 14058 -7178 14614
rect -6774 709082 -6218 709638
rect -6774 676338 -6218 676894
rect -6774 640338 -6218 640894
rect -6774 604338 -6218 604894
rect -6774 568338 -6218 568894
rect -6774 532338 -6218 532894
rect -6774 496338 -6218 496894
rect -6774 460338 -6218 460894
rect -6774 424338 -6218 424894
rect -6774 388338 -6218 388894
rect -6774 352338 -6218 352894
rect -6774 316338 -6218 316894
rect -6774 280338 -6218 280894
rect -6774 244338 -6218 244894
rect -6774 208338 -6218 208894
rect -6774 172338 -6218 172894
rect -6774 136338 -6218 136894
rect -6774 100338 -6218 100894
rect -6774 64338 -6218 64894
rect -6774 28338 -6218 28894
rect -5814 708122 -5258 708678
rect 9266 708122 9822 708678
rect -5814 694338 -5258 694894
rect -5814 658338 -5258 658894
rect -5814 622338 -5258 622894
rect -5814 586338 -5258 586894
rect -5814 550338 -5258 550894
rect -5814 514338 -5258 514894
rect -5814 478338 -5258 478894
rect -5814 442338 -5258 442894
rect -5814 406338 -5258 406894
rect -5814 370338 -5258 370894
rect -5814 334338 -5258 334894
rect -5814 298338 -5258 298894
rect -5814 262338 -5258 262894
rect -5814 226338 -5258 226894
rect -5814 190338 -5258 190894
rect -5814 154338 -5258 154894
rect -5814 118338 -5258 118894
rect -5814 82338 -5258 82894
rect -5814 46338 -5258 46894
rect -5814 10338 -5258 10894
rect -4854 707162 -4298 707718
rect -4854 672618 -4298 673174
rect -4854 636618 -4298 637174
rect -4854 600618 -4298 601174
rect -4854 564618 -4298 565174
rect -4854 528618 -4298 529174
rect -4854 492618 -4298 493174
rect -4854 456618 -4298 457174
rect -4854 420618 -4298 421174
rect -4854 384618 -4298 385174
rect -4854 348618 -4298 349174
rect -4854 312618 -4298 313174
rect -4854 276618 -4298 277174
rect -4854 240618 -4298 241174
rect -4854 204618 -4298 205174
rect -4854 168618 -4298 169174
rect -4854 132618 -4298 133174
rect -4854 96618 -4298 97174
rect -4854 60618 -4298 61174
rect -4854 24618 -4298 25174
rect -3894 706202 -3338 706758
rect 5546 706202 6102 706758
rect -3894 690618 -3338 691174
rect -3894 654618 -3338 655174
rect -3894 618618 -3338 619174
rect -3894 582618 -3338 583174
rect -3894 546618 -3338 547174
rect -3894 510618 -3338 511174
rect -3894 474618 -3338 475174
rect -3894 438618 -3338 439174
rect -3894 402618 -3338 403174
rect -3894 366618 -3338 367174
rect -3894 330618 -3338 331174
rect -3894 294618 -3338 295174
rect -3894 258618 -3338 259174
rect -3894 222618 -3338 223174
rect -3894 186618 -3338 187174
rect -3894 150618 -3338 151174
rect -3894 114618 -3338 115174
rect -3894 78618 -3338 79174
rect -3894 42618 -3338 43174
rect -3894 6618 -3338 7174
rect -2934 705242 -2378 705798
rect -2934 668898 -2378 669454
rect -2934 632898 -2378 633454
rect -2934 596898 -2378 597454
rect -2934 560898 -2378 561454
rect -2934 524898 -2378 525454
rect -2934 488898 -2378 489454
rect -2934 452898 -2378 453454
rect -2934 416898 -2378 417454
rect -2934 380898 -2378 381454
rect -2934 344898 -2378 345454
rect -2934 308898 -2378 309454
rect -2934 272898 -2378 273454
rect -2934 236898 -2378 237454
rect -2934 200898 -2378 201454
rect -2934 164898 -2378 165454
rect -2934 128898 -2378 129454
rect -2934 92898 -2378 93454
rect -2934 56898 -2378 57454
rect -2934 20898 -2378 21454
rect -1974 704282 -1418 704838
rect -1974 686898 -1418 687454
rect -1974 650898 -1418 651454
rect -1974 614898 -1418 615454
rect -1974 578898 -1418 579454
rect -1974 542898 -1418 543454
rect -1974 506898 -1418 507454
rect -1974 470898 -1418 471454
rect -1974 434898 -1418 435454
rect -1974 398898 -1418 399454
rect -1974 362898 -1418 363454
rect -1974 326898 -1418 327454
rect -1974 290898 -1418 291454
rect -1974 254898 -1418 255454
rect -1974 218898 -1418 219454
rect -1974 182898 -1418 183454
rect -1974 146898 -1418 147454
rect -1974 110898 -1418 111454
rect -1974 74898 -1418 75454
rect -1974 38898 -1418 39454
rect -1974 2898 -1418 3454
rect -1974 -902 -1418 -346
rect 1826 704282 2382 704838
rect 1826 686898 2382 687454
rect 1826 650898 2382 651454
rect 1826 614898 2382 615454
rect 1826 578898 2382 579454
rect 1826 542898 2382 543454
rect 1826 506898 2382 507454
rect 1826 470898 2382 471454
rect 1826 434898 2382 435454
rect 1826 398898 2382 399454
rect 1826 362898 2382 363454
rect 1826 326898 2382 327454
rect 1826 290898 2382 291454
rect 1826 254898 2382 255454
rect 1826 218898 2382 219454
rect 1826 182898 2382 183454
rect 1826 146898 2382 147454
rect 1826 110898 2382 111454
rect 1826 74898 2382 75454
rect 1826 38898 2382 39454
rect 1826 2898 2382 3454
rect 1826 -902 2382 -346
rect -2934 -1862 -2378 -1306
rect 5546 690618 6102 691174
rect 5546 654618 6102 655174
rect 5546 618618 6102 619174
rect 5546 582618 6102 583174
rect 5546 546618 6102 547174
rect 5546 510618 6102 511174
rect 5546 474618 6102 475174
rect 5546 438618 6102 439174
rect 5546 402618 6102 403174
rect 5546 366618 6102 367174
rect 5546 330618 6102 331174
rect 5546 294618 6102 295174
rect 5546 258618 6102 259174
rect 5546 222618 6102 223174
rect 5546 186618 6102 187174
rect 5546 150618 6102 151174
rect 5546 114618 6102 115174
rect 5546 78618 6102 79174
rect 5546 42618 6102 43174
rect 5546 6618 6102 7174
rect -3894 -2822 -3338 -2266
rect 5546 -2822 6102 -2266
rect -4854 -3782 -4298 -3226
rect 9266 694338 9822 694894
rect 9266 658338 9822 658894
rect 9266 622338 9822 622894
rect 9266 586338 9822 586894
rect 9266 550338 9822 550894
rect 9266 514338 9822 514894
rect 9266 478338 9822 478894
rect 9266 442338 9822 442894
rect 9266 406338 9822 406894
rect 9266 370338 9822 370894
rect 9266 334338 9822 334894
rect 9266 298338 9822 298894
rect 9266 262338 9822 262894
rect 9266 226338 9822 226894
rect 9266 190338 9822 190894
rect 9266 154338 9822 154894
rect 9266 118338 9822 118894
rect 9266 82338 9822 82894
rect 9266 46338 9822 46894
rect 9266 10338 9822 10894
rect -5814 -4742 -5258 -4186
rect 9266 -4742 9822 -4186
rect -6774 -5702 -6218 -5146
rect 30986 711002 31542 711558
rect 27266 709082 27822 709638
rect 23546 707162 24102 707718
rect 12986 698058 13542 698614
rect 12986 662058 13542 662614
rect 12986 626058 13542 626614
rect 12986 590058 13542 590614
rect 12986 554058 13542 554614
rect 12986 518058 13542 518614
rect 12986 482058 13542 482614
rect 12986 446058 13542 446614
rect 12986 410058 13542 410614
rect 12986 374058 13542 374614
rect 12986 338058 13542 338614
rect 12986 302058 13542 302614
rect 12986 266058 13542 266614
rect 12986 230058 13542 230614
rect 12986 194058 13542 194614
rect 12986 158058 13542 158614
rect 12986 122058 13542 122614
rect 12986 86058 13542 86614
rect 12986 50058 13542 50614
rect 12986 14058 13542 14614
rect -7734 -6662 -7178 -6106
rect 19826 705242 20382 705798
rect 19826 668898 20382 669454
rect 19826 632898 20382 633454
rect 19826 596898 20382 597454
rect 19826 560898 20382 561454
rect 19826 524898 20382 525454
rect 19826 488898 20382 489454
rect 19826 452898 20382 453454
rect 19826 416898 20382 417454
rect 19826 380898 20382 381454
rect 19826 344898 20382 345454
rect 19826 308898 20382 309454
rect 19826 272898 20382 273454
rect 19826 236898 20382 237454
rect 19826 200898 20382 201454
rect 19826 164898 20382 165454
rect 19826 128898 20382 129454
rect 19826 92898 20382 93454
rect 19826 56898 20382 57454
rect 19826 20898 20382 21454
rect 19826 -1862 20382 -1306
rect 23546 672618 24102 673174
rect 23546 636618 24102 637174
rect 23546 600618 24102 601174
rect 23546 564618 24102 565174
rect 23546 528618 24102 529174
rect 23546 492618 24102 493174
rect 23546 456618 24102 457174
rect 23546 420618 24102 421174
rect 23546 384618 24102 385174
rect 23546 348618 24102 349174
rect 23546 312618 24102 313174
rect 23546 276618 24102 277174
rect 23546 240618 24102 241174
rect 23546 204618 24102 205174
rect 23546 168618 24102 169174
rect 23546 132618 24102 133174
rect 23546 96618 24102 97174
rect 23546 60618 24102 61174
rect 23546 24618 24102 25174
rect 23546 -3782 24102 -3226
rect 27266 676338 27822 676894
rect 27266 640338 27822 640894
rect 27266 604338 27822 604894
rect 27266 568338 27822 568894
rect 27266 532338 27822 532894
rect 27266 496338 27822 496894
rect 27266 460338 27822 460894
rect 27266 424338 27822 424894
rect 27266 388338 27822 388894
rect 27266 352338 27822 352894
rect 27266 316338 27822 316894
rect 27266 280338 27822 280894
rect 27266 244338 27822 244894
rect 27266 208338 27822 208894
rect 27266 172338 27822 172894
rect 27266 136338 27822 136894
rect 27266 100338 27822 100894
rect 27266 64338 27822 64894
rect 27266 28338 27822 28894
rect 27266 -5702 27822 -5146
rect 48986 710042 49542 710598
rect 45266 708122 45822 708678
rect 41546 706202 42102 706758
rect 30986 680058 31542 680614
rect 30986 644058 31542 644614
rect 30986 608058 31542 608614
rect 30986 572058 31542 572614
rect 30986 536058 31542 536614
rect 30986 500058 31542 500614
rect 30986 464058 31542 464614
rect 30986 428058 31542 428614
rect 30986 392058 31542 392614
rect 30986 356058 31542 356614
rect 30986 320058 31542 320614
rect 30986 284058 31542 284614
rect 30986 248058 31542 248614
rect 30986 212058 31542 212614
rect 30986 176058 31542 176614
rect 30986 140058 31542 140614
rect 30986 104058 31542 104614
rect 30986 68058 31542 68614
rect 30986 32058 31542 32614
rect 12986 -6662 13542 -6106
rect -8694 -7622 -8138 -7066
rect 37826 704282 38382 704838
rect 37826 686898 38382 687454
rect 37826 650898 38382 651454
rect 37826 614898 38382 615454
rect 37826 578898 38382 579454
rect 37826 542898 38382 543454
rect 37826 506898 38382 507454
rect 37826 470898 38382 471454
rect 37826 434898 38382 435454
rect 37826 398898 38382 399454
rect 37826 362898 38382 363454
rect 37826 326898 38382 327454
rect 37826 290898 38382 291454
rect 37826 254898 38382 255454
rect 37826 218898 38382 219454
rect 37826 182898 38382 183454
rect 37826 146898 38382 147454
rect 37826 110898 38382 111454
rect 37826 74898 38382 75454
rect 37826 38898 38382 39454
rect 37826 2898 38382 3454
rect 37826 -902 38382 -346
rect 41546 690618 42102 691174
rect 41546 654618 42102 655174
rect 41546 618618 42102 619174
rect 41546 582618 42102 583174
rect 41546 546618 42102 547174
rect 41546 510618 42102 511174
rect 41546 474618 42102 475174
rect 41546 438618 42102 439174
rect 41546 402618 42102 403174
rect 41546 366618 42102 367174
rect 41546 330618 42102 331174
rect 41546 294618 42102 295174
rect 41546 258618 42102 259174
rect 41546 222618 42102 223174
rect 41546 186618 42102 187174
rect 41546 150618 42102 151174
rect 41546 114618 42102 115174
rect 41546 78618 42102 79174
rect 41546 42618 42102 43174
rect 41546 6618 42102 7174
rect 41546 -2822 42102 -2266
rect 45266 694338 45822 694894
rect 45266 658338 45822 658894
rect 45266 622338 45822 622894
rect 45266 586338 45822 586894
rect 45266 550338 45822 550894
rect 45266 514338 45822 514894
rect 45266 478338 45822 478894
rect 45266 442338 45822 442894
rect 45266 406338 45822 406894
rect 45266 370338 45822 370894
rect 45266 334338 45822 334894
rect 45266 298338 45822 298894
rect 45266 262338 45822 262894
rect 45266 226338 45822 226894
rect 45266 190338 45822 190894
rect 45266 154338 45822 154894
rect 45266 118338 45822 118894
rect 45266 82338 45822 82894
rect 45266 46338 45822 46894
rect 45266 10338 45822 10894
rect 45266 -4742 45822 -4186
rect 66986 711002 67542 711558
rect 63266 709082 63822 709638
rect 59546 707162 60102 707718
rect 48986 698058 49542 698614
rect 48986 662058 49542 662614
rect 48986 626058 49542 626614
rect 48986 590058 49542 590614
rect 48986 554058 49542 554614
rect 48986 518058 49542 518614
rect 48986 482058 49542 482614
rect 48986 446058 49542 446614
rect 48986 410058 49542 410614
rect 48986 374058 49542 374614
rect 48986 338058 49542 338614
rect 48986 302058 49542 302614
rect 48986 266058 49542 266614
rect 48986 230058 49542 230614
rect 48986 194058 49542 194614
rect 48986 158058 49542 158614
rect 48986 122058 49542 122614
rect 48986 86058 49542 86614
rect 48986 50058 49542 50614
rect 48986 14058 49542 14614
rect 30986 -7622 31542 -7066
rect 55826 705242 56382 705798
rect 55826 668898 56382 669454
rect 55826 632898 56382 633454
rect 55826 596898 56382 597454
rect 55826 560898 56382 561454
rect 55826 524898 56382 525454
rect 55826 488898 56382 489454
rect 55826 452898 56382 453454
rect 55826 416898 56382 417454
rect 55826 380898 56382 381454
rect 55826 344898 56382 345454
rect 55826 308898 56382 309454
rect 55826 272898 56382 273454
rect 55826 236898 56382 237454
rect 55826 200898 56382 201454
rect 55826 164898 56382 165454
rect 55826 128898 56382 129454
rect 55826 92898 56382 93454
rect 55826 56898 56382 57454
rect 55826 20898 56382 21454
rect 55826 -1862 56382 -1306
rect 59546 672618 60102 673174
rect 59546 636618 60102 637174
rect 59546 600618 60102 601174
rect 59546 564618 60102 565174
rect 59546 528618 60102 529174
rect 59546 492618 60102 493174
rect 59546 456618 60102 457174
rect 59546 420618 60102 421174
rect 59546 384618 60102 385174
rect 59546 348618 60102 349174
rect 59546 312618 60102 313174
rect 59546 276618 60102 277174
rect 59546 240618 60102 241174
rect 59546 204618 60102 205174
rect 59546 168618 60102 169174
rect 59546 132618 60102 133174
rect 59546 96618 60102 97174
rect 59546 60618 60102 61174
rect 59546 24618 60102 25174
rect 59546 -3782 60102 -3226
rect 63266 676338 63822 676894
rect 63266 640338 63822 640894
rect 63266 604338 63822 604894
rect 63266 568338 63822 568894
rect 63266 532338 63822 532894
rect 63266 496338 63822 496894
rect 63266 460338 63822 460894
rect 63266 424338 63822 424894
rect 63266 388338 63822 388894
rect 63266 352338 63822 352894
rect 63266 316338 63822 316894
rect 63266 280338 63822 280894
rect 63266 244338 63822 244894
rect 63266 208338 63822 208894
rect 63266 172338 63822 172894
rect 63266 136338 63822 136894
rect 63266 100338 63822 100894
rect 63266 64338 63822 64894
rect 63266 28338 63822 28894
rect 63266 -5702 63822 -5146
rect 84986 710042 85542 710598
rect 81266 708122 81822 708678
rect 77546 706202 78102 706758
rect 66986 680058 67542 680614
rect 66986 644058 67542 644614
rect 66986 608058 67542 608614
rect 66986 572058 67542 572614
rect 66986 536058 67542 536614
rect 66986 500058 67542 500614
rect 66986 464058 67542 464614
rect 66986 428058 67542 428614
rect 66986 392058 67542 392614
rect 66986 356058 67542 356614
rect 66986 320058 67542 320614
rect 66986 284058 67542 284614
rect 66986 248058 67542 248614
rect 66986 212058 67542 212614
rect 66986 176058 67542 176614
rect 66986 140058 67542 140614
rect 66986 104058 67542 104614
rect 66986 68058 67542 68614
rect 66986 32058 67542 32614
rect 48986 -6662 49542 -6106
rect 73826 704282 74382 704838
rect 73826 686898 74382 687454
rect 73826 650898 74382 651454
rect 73826 614898 74382 615454
rect 73826 578898 74382 579454
rect 73826 542898 74382 543454
rect 73826 506898 74382 507454
rect 73826 470898 74382 471454
rect 73826 434898 74382 435454
rect 73826 398898 74382 399454
rect 73826 362898 74382 363454
rect 73826 326898 74382 327454
rect 73826 290898 74382 291454
rect 73826 254898 74382 255454
rect 73826 218898 74382 219454
rect 73826 182898 74382 183454
rect 73826 146898 74382 147454
rect 73826 110898 74382 111454
rect 73826 74898 74382 75454
rect 73826 38898 74382 39454
rect 73826 2898 74382 3454
rect 73826 -902 74382 -346
rect 77546 690618 78102 691174
rect 77546 654618 78102 655174
rect 77546 618618 78102 619174
rect 77546 582618 78102 583174
rect 77546 546618 78102 547174
rect 77546 510618 78102 511174
rect 77546 474618 78102 475174
rect 77546 438618 78102 439174
rect 77546 402618 78102 403174
rect 77546 366618 78102 367174
rect 77546 330618 78102 331174
rect 77546 294618 78102 295174
rect 77546 258618 78102 259174
rect 77546 222618 78102 223174
rect 77546 186618 78102 187174
rect 77546 150618 78102 151174
rect 77546 114618 78102 115174
rect 77546 78618 78102 79174
rect 77546 42618 78102 43174
rect 77546 6618 78102 7174
rect 77546 -2822 78102 -2266
rect 81266 694338 81822 694894
rect 81266 658338 81822 658894
rect 81266 622338 81822 622894
rect 81266 586338 81822 586894
rect 81266 550338 81822 550894
rect 81266 514338 81822 514894
rect 81266 478338 81822 478894
rect 81266 442338 81822 442894
rect 81266 406338 81822 406894
rect 81266 370338 81822 370894
rect 81266 334338 81822 334894
rect 81266 298338 81822 298894
rect 81266 262338 81822 262894
rect 81266 226338 81822 226894
rect 81266 190338 81822 190894
rect 81266 154338 81822 154894
rect 81266 118338 81822 118894
rect 81266 82338 81822 82894
rect 81266 46338 81822 46894
rect 81266 10338 81822 10894
rect 81266 -4742 81822 -4186
rect 102986 711002 103542 711558
rect 99266 709082 99822 709638
rect 95546 707162 96102 707718
rect 84986 698058 85542 698614
rect 84986 662058 85542 662614
rect 84986 626058 85542 626614
rect 84986 590058 85542 590614
rect 84986 554058 85542 554614
rect 84986 518058 85542 518614
rect 84986 482058 85542 482614
rect 84986 446058 85542 446614
rect 84986 410058 85542 410614
rect 84986 374058 85542 374614
rect 84986 338058 85542 338614
rect 84986 302058 85542 302614
rect 84986 266058 85542 266614
rect 84986 230058 85542 230614
rect 84986 194058 85542 194614
rect 84986 158058 85542 158614
rect 84986 122058 85542 122614
rect 84986 86058 85542 86614
rect 84986 50058 85542 50614
rect 84986 14058 85542 14614
rect 66986 -7622 67542 -7066
rect 91826 705242 92382 705798
rect 91826 668898 92382 669454
rect 91826 632898 92382 633454
rect 91826 596898 92382 597454
rect 91826 560898 92382 561454
rect 91826 524898 92382 525454
rect 91826 488898 92382 489454
rect 91826 452898 92382 453454
rect 91826 416898 92382 417454
rect 91826 380898 92382 381454
rect 91826 344898 92382 345454
rect 91826 308898 92382 309454
rect 91826 272898 92382 273454
rect 91826 236898 92382 237454
rect 91826 200898 92382 201454
rect 91826 164898 92382 165454
rect 91826 128898 92382 129454
rect 91826 92898 92382 93454
rect 91826 56898 92382 57454
rect 91826 20898 92382 21454
rect 91826 -1862 92382 -1306
rect 95546 672618 96102 673174
rect 95546 636618 96102 637174
rect 95546 600618 96102 601174
rect 95546 564618 96102 565174
rect 95546 528618 96102 529174
rect 95546 492618 96102 493174
rect 95546 456618 96102 457174
rect 95546 420618 96102 421174
rect 95546 384618 96102 385174
rect 95546 348618 96102 349174
rect 95546 312618 96102 313174
rect 95546 276618 96102 277174
rect 95546 240618 96102 241174
rect 95546 204618 96102 205174
rect 95546 168618 96102 169174
rect 95546 132618 96102 133174
rect 95546 96618 96102 97174
rect 95546 60618 96102 61174
rect 95546 24618 96102 25174
rect 95546 -3782 96102 -3226
rect 99266 676338 99822 676894
rect 99266 640338 99822 640894
rect 99266 604338 99822 604894
rect 99266 568338 99822 568894
rect 99266 532338 99822 532894
rect 99266 496338 99822 496894
rect 99266 460338 99822 460894
rect 99266 424338 99822 424894
rect 99266 388338 99822 388894
rect 99266 352338 99822 352894
rect 99266 316338 99822 316894
rect 99266 280338 99822 280894
rect 99266 244338 99822 244894
rect 99266 208338 99822 208894
rect 99266 172338 99822 172894
rect 99266 136338 99822 136894
rect 99266 100338 99822 100894
rect 99266 64338 99822 64894
rect 99266 28338 99822 28894
rect 99266 -5702 99822 -5146
rect 120986 710042 121542 710598
rect 117266 708122 117822 708678
rect 113546 706202 114102 706758
rect 102986 680058 103542 680614
rect 102986 644058 103542 644614
rect 102986 608058 103542 608614
rect 102986 572058 103542 572614
rect 102986 536058 103542 536614
rect 102986 500058 103542 500614
rect 102986 464058 103542 464614
rect 102986 428058 103542 428614
rect 102986 392058 103542 392614
rect 102986 356058 103542 356614
rect 102986 320058 103542 320614
rect 102986 284058 103542 284614
rect 102986 248058 103542 248614
rect 102986 212058 103542 212614
rect 102986 176058 103542 176614
rect 102986 140058 103542 140614
rect 102986 104058 103542 104614
rect 102986 68058 103542 68614
rect 102986 32058 103542 32614
rect 84986 -6662 85542 -6106
rect 109826 704282 110382 704838
rect 109826 686898 110382 687454
rect 109826 650898 110382 651454
rect 109826 614898 110382 615454
rect 109826 578898 110382 579454
rect 109826 542898 110382 543454
rect 109826 506898 110382 507454
rect 109826 470898 110382 471454
rect 109826 434898 110382 435454
rect 109826 398898 110382 399454
rect 109826 362898 110382 363454
rect 109826 326898 110382 327454
rect 109826 290898 110382 291454
rect 109826 254898 110382 255454
rect 109826 218898 110382 219454
rect 109826 182898 110382 183454
rect 109826 146898 110382 147454
rect 109826 110898 110382 111454
rect 109826 74898 110382 75454
rect 109826 38898 110382 39454
rect 109826 2898 110382 3454
rect 109826 -902 110382 -346
rect 113546 690618 114102 691174
rect 113546 654618 114102 655174
rect 113546 618618 114102 619174
rect 113546 582618 114102 583174
rect 113546 546618 114102 547174
rect 113546 510618 114102 511174
rect 113546 474618 114102 475174
rect 113546 438618 114102 439174
rect 113546 402618 114102 403174
rect 113546 366618 114102 367174
rect 113546 330618 114102 331174
rect 113546 294618 114102 295174
rect 113546 258618 114102 259174
rect 113546 222618 114102 223174
rect 113546 186618 114102 187174
rect 113546 150618 114102 151174
rect 113546 114618 114102 115174
rect 113546 78618 114102 79174
rect 113546 42618 114102 43174
rect 113546 6618 114102 7174
rect 113546 -2822 114102 -2266
rect 117266 694338 117822 694894
rect 117266 658338 117822 658894
rect 117266 622338 117822 622894
rect 117266 586338 117822 586894
rect 117266 550338 117822 550894
rect 117266 514338 117822 514894
rect 117266 478338 117822 478894
rect 117266 442338 117822 442894
rect 117266 406338 117822 406894
rect 117266 370338 117822 370894
rect 117266 334338 117822 334894
rect 117266 298338 117822 298894
rect 117266 262338 117822 262894
rect 117266 226338 117822 226894
rect 117266 190338 117822 190894
rect 117266 154338 117822 154894
rect 117266 118338 117822 118894
rect 117266 82338 117822 82894
rect 117266 46338 117822 46894
rect 117266 10338 117822 10894
rect 117266 -4742 117822 -4186
rect 138986 711002 139542 711558
rect 135266 709082 135822 709638
rect 131546 707162 132102 707718
rect 120986 698058 121542 698614
rect 120986 662058 121542 662614
rect 120986 626058 121542 626614
rect 120986 590058 121542 590614
rect 120986 554058 121542 554614
rect 120986 518058 121542 518614
rect 120986 482058 121542 482614
rect 120986 446058 121542 446614
rect 120986 410058 121542 410614
rect 120986 374058 121542 374614
rect 120986 338058 121542 338614
rect 120986 302058 121542 302614
rect 120986 266058 121542 266614
rect 120986 230058 121542 230614
rect 120986 194058 121542 194614
rect 120986 158058 121542 158614
rect 120986 122058 121542 122614
rect 120986 86058 121542 86614
rect 120986 50058 121542 50614
rect 120986 14058 121542 14614
rect 102986 -7622 103542 -7066
rect 127826 705242 128382 705798
rect 127826 668898 128382 669454
rect 127826 632898 128382 633454
rect 127826 596898 128382 597454
rect 127826 560898 128382 561454
rect 127826 524898 128382 525454
rect 127826 488898 128382 489454
rect 127826 452898 128382 453454
rect 127826 416898 128382 417454
rect 127826 380898 128382 381454
rect 127826 344898 128382 345454
rect 127826 308898 128382 309454
rect 127826 272898 128382 273454
rect 127826 236898 128382 237454
rect 127826 200898 128382 201454
rect 127826 164898 128382 165454
rect 127826 128898 128382 129454
rect 127826 92898 128382 93454
rect 127826 56898 128382 57454
rect 127826 20898 128382 21454
rect 127826 -1862 128382 -1306
rect 131546 672618 132102 673174
rect 131546 636618 132102 637174
rect 131546 600618 132102 601174
rect 131546 564618 132102 565174
rect 131546 528618 132102 529174
rect 131546 492618 132102 493174
rect 131546 456618 132102 457174
rect 131546 420618 132102 421174
rect 131546 384618 132102 385174
rect 131546 348618 132102 349174
rect 131546 312618 132102 313174
rect 131546 276618 132102 277174
rect 131546 240618 132102 241174
rect 131546 204618 132102 205174
rect 131546 168618 132102 169174
rect 131546 132618 132102 133174
rect 131546 96618 132102 97174
rect 131546 60618 132102 61174
rect 131546 24618 132102 25174
rect 131546 -3782 132102 -3226
rect 135266 676338 135822 676894
rect 135266 640338 135822 640894
rect 135266 604338 135822 604894
rect 135266 568338 135822 568894
rect 135266 532338 135822 532894
rect 135266 496338 135822 496894
rect 135266 460338 135822 460894
rect 135266 424338 135822 424894
rect 135266 388338 135822 388894
rect 135266 352338 135822 352894
rect 135266 316338 135822 316894
rect 135266 280338 135822 280894
rect 135266 244338 135822 244894
rect 135266 208338 135822 208894
rect 135266 172338 135822 172894
rect 135266 136338 135822 136894
rect 135266 100338 135822 100894
rect 135266 64338 135822 64894
rect 135266 28338 135822 28894
rect 135266 -5702 135822 -5146
rect 156986 710042 157542 710598
rect 153266 708122 153822 708678
rect 149546 706202 150102 706758
rect 138986 680058 139542 680614
rect 138986 644058 139542 644614
rect 138986 608058 139542 608614
rect 138986 572058 139542 572614
rect 138986 536058 139542 536614
rect 138986 500058 139542 500614
rect 138986 464058 139542 464614
rect 138986 428058 139542 428614
rect 138986 392058 139542 392614
rect 138986 356058 139542 356614
rect 138986 320058 139542 320614
rect 138986 284058 139542 284614
rect 138986 248058 139542 248614
rect 138986 212058 139542 212614
rect 138986 176058 139542 176614
rect 138986 140058 139542 140614
rect 138986 104058 139542 104614
rect 138986 68058 139542 68614
rect 138986 32058 139542 32614
rect 120986 -6662 121542 -6106
rect 145826 704282 146382 704838
rect 145826 686898 146382 687454
rect 145826 650898 146382 651454
rect 145826 614898 146382 615454
rect 145826 578898 146382 579454
rect 145826 542898 146382 543454
rect 145826 506898 146382 507454
rect 145826 470898 146382 471454
rect 145826 434898 146382 435454
rect 145826 398898 146382 399454
rect 145826 362898 146382 363454
rect 145826 326898 146382 327454
rect 145826 290898 146382 291454
rect 145826 254898 146382 255454
rect 145826 218898 146382 219454
rect 145826 182898 146382 183454
rect 145826 146898 146382 147454
rect 145826 110898 146382 111454
rect 145826 74898 146382 75454
rect 145826 38898 146382 39454
rect 145826 2898 146382 3454
rect 145826 -902 146382 -346
rect 149546 690618 150102 691174
rect 149546 654618 150102 655174
rect 149546 618618 150102 619174
rect 149546 582618 150102 583174
rect 149546 546618 150102 547174
rect 149546 510618 150102 511174
rect 149546 474618 150102 475174
rect 149546 438618 150102 439174
rect 149546 402618 150102 403174
rect 149546 366618 150102 367174
rect 149546 330618 150102 331174
rect 149546 294618 150102 295174
rect 149546 258618 150102 259174
rect 149546 222618 150102 223174
rect 149546 186618 150102 187174
rect 149546 150618 150102 151174
rect 149546 114618 150102 115174
rect 149546 78618 150102 79174
rect 149546 42618 150102 43174
rect 149546 6618 150102 7174
rect 149546 -2822 150102 -2266
rect 153266 694338 153822 694894
rect 153266 658338 153822 658894
rect 153266 622338 153822 622894
rect 153266 586338 153822 586894
rect 153266 550338 153822 550894
rect 153266 514338 153822 514894
rect 153266 478338 153822 478894
rect 153266 442338 153822 442894
rect 153266 406338 153822 406894
rect 153266 370338 153822 370894
rect 153266 334338 153822 334894
rect 153266 298338 153822 298894
rect 153266 262338 153822 262894
rect 153266 226338 153822 226894
rect 153266 190338 153822 190894
rect 153266 154338 153822 154894
rect 153266 118338 153822 118894
rect 153266 82338 153822 82894
rect 153266 46338 153822 46894
rect 153266 10338 153822 10894
rect 153266 -4742 153822 -4186
rect 174986 711002 175542 711558
rect 171266 709082 171822 709638
rect 167546 707162 168102 707718
rect 156986 698058 157542 698614
rect 156986 662058 157542 662614
rect 156986 626058 157542 626614
rect 156986 590058 157542 590614
rect 156986 554058 157542 554614
rect 156986 518058 157542 518614
rect 156986 482058 157542 482614
rect 156986 446058 157542 446614
rect 156986 410058 157542 410614
rect 156986 374058 157542 374614
rect 156986 338058 157542 338614
rect 156986 302058 157542 302614
rect 156986 266058 157542 266614
rect 156986 230058 157542 230614
rect 156986 194058 157542 194614
rect 156986 158058 157542 158614
rect 156986 122058 157542 122614
rect 156986 86058 157542 86614
rect 156986 50058 157542 50614
rect 156986 14058 157542 14614
rect 138986 -7622 139542 -7066
rect 163826 705242 164382 705798
rect 163826 668898 164382 669454
rect 163826 632898 164382 633454
rect 163826 596898 164382 597454
rect 163826 560898 164382 561454
rect 163826 524898 164382 525454
rect 163826 488898 164382 489454
rect 163826 452898 164382 453454
rect 163826 416898 164382 417454
rect 163826 380898 164382 381454
rect 163826 344898 164382 345454
rect 163826 308898 164382 309454
rect 163826 272898 164382 273454
rect 163826 236898 164382 237454
rect 163826 200898 164382 201454
rect 163826 164898 164382 165454
rect 163826 128898 164382 129454
rect 163826 92898 164382 93454
rect 163826 56898 164382 57454
rect 163826 20898 164382 21454
rect 163826 -1862 164382 -1306
rect 167546 672618 168102 673174
rect 167546 636618 168102 637174
rect 167546 600618 168102 601174
rect 167546 564618 168102 565174
rect 167546 528618 168102 529174
rect 167546 492618 168102 493174
rect 167546 456618 168102 457174
rect 167546 420618 168102 421174
rect 167546 384618 168102 385174
rect 167546 348618 168102 349174
rect 167546 312618 168102 313174
rect 167546 276618 168102 277174
rect 167546 240618 168102 241174
rect 167546 204618 168102 205174
rect 167546 168618 168102 169174
rect 167546 132618 168102 133174
rect 167546 96618 168102 97174
rect 167546 60618 168102 61174
rect 167546 24618 168102 25174
rect 167546 -3782 168102 -3226
rect 171266 676338 171822 676894
rect 171266 640338 171822 640894
rect 171266 604338 171822 604894
rect 171266 568338 171822 568894
rect 171266 532338 171822 532894
rect 171266 496338 171822 496894
rect 171266 460338 171822 460894
rect 171266 424338 171822 424894
rect 171266 388338 171822 388894
rect 171266 352338 171822 352894
rect 171266 316338 171822 316894
rect 171266 280338 171822 280894
rect 171266 244338 171822 244894
rect 171266 208338 171822 208894
rect 171266 172338 171822 172894
rect 171266 136338 171822 136894
rect 171266 100338 171822 100894
rect 171266 64338 171822 64894
rect 171266 28338 171822 28894
rect 171266 -5702 171822 -5146
rect 192986 710042 193542 710598
rect 189266 708122 189822 708678
rect 185546 706202 186102 706758
rect 174986 680058 175542 680614
rect 174986 644058 175542 644614
rect 174986 608058 175542 608614
rect 174986 572058 175542 572614
rect 174986 536058 175542 536614
rect 174986 500058 175542 500614
rect 174986 464058 175542 464614
rect 174986 428058 175542 428614
rect 174986 392058 175542 392614
rect 174986 356058 175542 356614
rect 174986 320058 175542 320614
rect 174986 284058 175542 284614
rect 174986 248058 175542 248614
rect 174986 212058 175542 212614
rect 174986 176058 175542 176614
rect 174986 140058 175542 140614
rect 174986 104058 175542 104614
rect 174986 68058 175542 68614
rect 174986 32058 175542 32614
rect 156986 -6662 157542 -6106
rect 181826 704282 182382 704838
rect 181826 686898 182382 687454
rect 181826 650898 182382 651454
rect 181826 614898 182382 615454
rect 181826 578898 182382 579454
rect 181826 542898 182382 543454
rect 181826 506898 182382 507454
rect 181826 470898 182382 471454
rect 181826 434898 182382 435454
rect 181826 398898 182382 399454
rect 181826 362898 182382 363454
rect 181826 326898 182382 327454
rect 181826 290898 182382 291454
rect 181826 254898 182382 255454
rect 181826 218898 182382 219454
rect 181826 182898 182382 183454
rect 181826 146898 182382 147454
rect 181826 110898 182382 111454
rect 181826 74898 182382 75454
rect 181826 38898 182382 39454
rect 181826 2898 182382 3454
rect 181826 -902 182382 -346
rect 185546 690618 186102 691174
rect 185546 654618 186102 655174
rect 185546 618618 186102 619174
rect 185546 582618 186102 583174
rect 185546 546618 186102 547174
rect 185546 510618 186102 511174
rect 185546 474618 186102 475174
rect 185546 438618 186102 439174
rect 185546 402618 186102 403174
rect 185546 366618 186102 367174
rect 185546 330618 186102 331174
rect 185546 294618 186102 295174
rect 185546 258618 186102 259174
rect 185546 222618 186102 223174
rect 185546 186618 186102 187174
rect 185546 150618 186102 151174
rect 185546 114618 186102 115174
rect 185546 78618 186102 79174
rect 185546 42618 186102 43174
rect 185546 6618 186102 7174
rect 185546 -2822 186102 -2266
rect 189266 694338 189822 694894
rect 189266 658338 189822 658894
rect 189266 622338 189822 622894
rect 189266 586338 189822 586894
rect 189266 550338 189822 550894
rect 189266 514338 189822 514894
rect 189266 478338 189822 478894
rect 189266 442338 189822 442894
rect 189266 406338 189822 406894
rect 189266 370338 189822 370894
rect 189266 334338 189822 334894
rect 189266 298338 189822 298894
rect 189266 262338 189822 262894
rect 189266 226338 189822 226894
rect 189266 190338 189822 190894
rect 189266 154338 189822 154894
rect 189266 118338 189822 118894
rect 189266 82338 189822 82894
rect 189266 46338 189822 46894
rect 189266 10338 189822 10894
rect 189266 -4742 189822 -4186
rect 210986 711002 211542 711558
rect 207266 709082 207822 709638
rect 203546 707162 204102 707718
rect 192986 698058 193542 698614
rect 192986 662058 193542 662614
rect 192986 626058 193542 626614
rect 192986 590058 193542 590614
rect 192986 554058 193542 554614
rect 192986 518058 193542 518614
rect 192986 482058 193542 482614
rect 192986 446058 193542 446614
rect 192986 410058 193542 410614
rect 192986 374058 193542 374614
rect 192986 338058 193542 338614
rect 192986 302058 193542 302614
rect 192986 266058 193542 266614
rect 192986 230058 193542 230614
rect 192986 194058 193542 194614
rect 192986 158058 193542 158614
rect 192986 122058 193542 122614
rect 192986 86058 193542 86614
rect 192986 50058 193542 50614
rect 192986 14058 193542 14614
rect 174986 -7622 175542 -7066
rect 199826 705242 200382 705798
rect 199826 668898 200382 669454
rect 199826 632898 200382 633454
rect 199826 596898 200382 597454
rect 199826 560898 200382 561454
rect 199826 524898 200382 525454
rect 199826 488898 200382 489454
rect 199826 452898 200382 453454
rect 199826 416898 200382 417454
rect 199826 380898 200382 381454
rect 199826 344898 200382 345454
rect 199826 308898 200382 309454
rect 199826 272898 200382 273454
rect 199826 236898 200382 237454
rect 199826 200898 200382 201454
rect 199826 164898 200382 165454
rect 199826 128898 200382 129454
rect 199826 92898 200382 93454
rect 199826 56898 200382 57454
rect 199826 20898 200382 21454
rect 199826 -1862 200382 -1306
rect 203546 672618 204102 673174
rect 203546 636618 204102 637174
rect 203546 600618 204102 601174
rect 203546 564618 204102 565174
rect 203546 528618 204102 529174
rect 203546 492618 204102 493174
rect 203546 456618 204102 457174
rect 203546 420618 204102 421174
rect 203546 384618 204102 385174
rect 203546 348618 204102 349174
rect 203546 312618 204102 313174
rect 203546 276618 204102 277174
rect 203546 240618 204102 241174
rect 203546 204618 204102 205174
rect 203546 168618 204102 169174
rect 203546 132618 204102 133174
rect 203546 96618 204102 97174
rect 203546 60618 204102 61174
rect 203546 24618 204102 25174
rect 203546 -3782 204102 -3226
rect 207266 676338 207822 676894
rect 207266 640338 207822 640894
rect 207266 604338 207822 604894
rect 207266 568338 207822 568894
rect 207266 532338 207822 532894
rect 207266 496338 207822 496894
rect 207266 460338 207822 460894
rect 207266 424338 207822 424894
rect 207266 388338 207822 388894
rect 207266 352338 207822 352894
rect 207266 316338 207822 316894
rect 207266 280338 207822 280894
rect 207266 244338 207822 244894
rect 207266 208338 207822 208894
rect 207266 172338 207822 172894
rect 207266 136338 207822 136894
rect 207266 100338 207822 100894
rect 207266 64338 207822 64894
rect 207266 28338 207822 28894
rect 207266 -5702 207822 -5146
rect 228986 710042 229542 710598
rect 225266 708122 225822 708678
rect 221546 706202 222102 706758
rect 210986 680058 211542 680614
rect 210986 644058 211542 644614
rect 210986 608058 211542 608614
rect 210986 572058 211542 572614
rect 210986 536058 211542 536614
rect 210986 500058 211542 500614
rect 210986 464058 211542 464614
rect 210986 428058 211542 428614
rect 210986 392058 211542 392614
rect 210986 356058 211542 356614
rect 210986 320058 211542 320614
rect 210986 284058 211542 284614
rect 210986 248058 211542 248614
rect 210986 212058 211542 212614
rect 210986 176058 211542 176614
rect 210986 140058 211542 140614
rect 210986 104058 211542 104614
rect 210986 68058 211542 68614
rect 210986 32058 211542 32614
rect 192986 -6662 193542 -6106
rect 217826 704282 218382 704838
rect 217826 686898 218382 687454
rect 217826 650898 218382 651454
rect 217826 614898 218382 615454
rect 217826 578898 218382 579454
rect 217826 542898 218382 543454
rect 217826 506898 218382 507454
rect 217826 470898 218382 471454
rect 217826 434898 218382 435454
rect 217826 398898 218382 399454
rect 217826 362898 218382 363454
rect 217826 326898 218382 327454
rect 217826 290898 218382 291454
rect 217826 254898 218382 255454
rect 217826 218898 218382 219454
rect 217826 182898 218382 183454
rect 217826 146898 218382 147454
rect 217826 110898 218382 111454
rect 217826 74898 218382 75454
rect 217826 38898 218382 39454
rect 217826 2898 218382 3454
rect 217826 -902 218382 -346
rect 221546 690618 222102 691174
rect 221546 654618 222102 655174
rect 221546 618618 222102 619174
rect 221546 582618 222102 583174
rect 221546 546618 222102 547174
rect 221546 510618 222102 511174
rect 221546 474618 222102 475174
rect 221546 438618 222102 439174
rect 221546 402618 222102 403174
rect 221546 366618 222102 367174
rect 221546 330618 222102 331174
rect 221546 294618 222102 295174
rect 221546 258618 222102 259174
rect 221546 222618 222102 223174
rect 221546 186618 222102 187174
rect 221546 150618 222102 151174
rect 221546 114618 222102 115174
rect 221546 78618 222102 79174
rect 221546 42618 222102 43174
rect 221546 6618 222102 7174
rect 221546 -2822 222102 -2266
rect 225266 694338 225822 694894
rect 225266 658338 225822 658894
rect 225266 622338 225822 622894
rect 225266 586338 225822 586894
rect 225266 550338 225822 550894
rect 225266 514338 225822 514894
rect 225266 478338 225822 478894
rect 225266 442338 225822 442894
rect 225266 406338 225822 406894
rect 225266 370338 225822 370894
rect 225266 334338 225822 334894
rect 225266 298338 225822 298894
rect 225266 262338 225822 262894
rect 225266 226338 225822 226894
rect 225266 190338 225822 190894
rect 225266 154338 225822 154894
rect 225266 118338 225822 118894
rect 225266 82338 225822 82894
rect 225266 46338 225822 46894
rect 225266 10338 225822 10894
rect 225266 -4742 225822 -4186
rect 246986 711002 247542 711558
rect 243266 709082 243822 709638
rect 239546 707162 240102 707718
rect 228986 698058 229542 698614
rect 228986 662058 229542 662614
rect 228986 626058 229542 626614
rect 228986 590058 229542 590614
rect 228986 554058 229542 554614
rect 228986 518058 229542 518614
rect 228986 482058 229542 482614
rect 228986 446058 229542 446614
rect 228986 410058 229542 410614
rect 235826 705242 236382 705798
rect 235826 668898 236382 669454
rect 235826 632898 236382 633454
rect 235826 596898 236382 597454
rect 235826 560898 236382 561454
rect 235826 524898 236382 525454
rect 235826 488898 236382 489454
rect 235826 452898 236382 453454
rect 235826 416898 236382 417454
rect 235826 380898 236382 381454
rect 239546 672618 240102 673174
rect 239546 636618 240102 637174
rect 239546 600618 240102 601174
rect 239546 564618 240102 565174
rect 239546 528618 240102 529174
rect 239546 492618 240102 493174
rect 239546 456618 240102 457174
rect 239546 420618 240102 421174
rect 239546 384618 240102 385174
rect 243266 676338 243822 676894
rect 243266 640338 243822 640894
rect 243266 604338 243822 604894
rect 243266 568338 243822 568894
rect 243266 532338 243822 532894
rect 243266 496338 243822 496894
rect 243266 460338 243822 460894
rect 243266 424338 243822 424894
rect 243266 388338 243822 388894
rect 264986 710042 265542 710598
rect 261266 708122 261822 708678
rect 257546 706202 258102 706758
rect 246986 680058 247542 680614
rect 246986 644058 247542 644614
rect 246986 608058 247542 608614
rect 246986 572058 247542 572614
rect 246986 536058 247542 536614
rect 246986 500058 247542 500614
rect 246986 464058 247542 464614
rect 246986 428058 247542 428614
rect 246986 392058 247542 392614
rect 253826 704282 254382 704838
rect 253826 686898 254382 687454
rect 253826 650898 254382 651454
rect 253826 614898 254382 615454
rect 253826 578898 254382 579454
rect 253826 542898 254382 543454
rect 253826 506898 254382 507454
rect 253826 470898 254382 471454
rect 253826 434898 254382 435454
rect 253826 398898 254382 399454
rect 257546 690618 258102 691174
rect 257546 654618 258102 655174
rect 257546 618618 258102 619174
rect 257546 582618 258102 583174
rect 257546 546618 258102 547174
rect 257546 510618 258102 511174
rect 257546 474618 258102 475174
rect 257546 438618 258102 439174
rect 257546 402618 258102 403174
rect 261266 694338 261822 694894
rect 261266 658338 261822 658894
rect 261266 622338 261822 622894
rect 261266 586338 261822 586894
rect 261266 550338 261822 550894
rect 261266 514338 261822 514894
rect 261266 478338 261822 478894
rect 261266 442338 261822 442894
rect 261266 406338 261822 406894
rect 282986 711002 283542 711558
rect 279266 709082 279822 709638
rect 275546 707162 276102 707718
rect 264986 698058 265542 698614
rect 264986 662058 265542 662614
rect 264986 626058 265542 626614
rect 264986 590058 265542 590614
rect 264986 554058 265542 554614
rect 264986 518058 265542 518614
rect 264986 482058 265542 482614
rect 264986 446058 265542 446614
rect 264986 410058 265542 410614
rect 271826 705242 272382 705798
rect 271826 668898 272382 669454
rect 271826 632898 272382 633454
rect 271826 596898 272382 597454
rect 271826 560898 272382 561454
rect 271826 524898 272382 525454
rect 271826 488898 272382 489454
rect 271826 452898 272382 453454
rect 271826 416898 272382 417454
rect 271826 380898 272382 381454
rect 275546 672618 276102 673174
rect 275546 636618 276102 637174
rect 275546 600618 276102 601174
rect 275546 564618 276102 565174
rect 275546 528618 276102 529174
rect 275546 492618 276102 493174
rect 275546 456618 276102 457174
rect 275546 420618 276102 421174
rect 275546 384618 276102 385174
rect 279266 676338 279822 676894
rect 279266 640338 279822 640894
rect 279266 604338 279822 604894
rect 279266 568338 279822 568894
rect 279266 532338 279822 532894
rect 279266 496338 279822 496894
rect 279266 460338 279822 460894
rect 279266 424338 279822 424894
rect 279266 388338 279822 388894
rect 300986 710042 301542 710598
rect 297266 708122 297822 708678
rect 293546 706202 294102 706758
rect 282986 680058 283542 680614
rect 282986 644058 283542 644614
rect 282986 608058 283542 608614
rect 282986 572058 283542 572614
rect 282986 536058 283542 536614
rect 282986 500058 283542 500614
rect 282986 464058 283542 464614
rect 282986 428058 283542 428614
rect 282986 392058 283542 392614
rect 289826 704282 290382 704838
rect 289826 686898 290382 687454
rect 289826 650898 290382 651454
rect 289826 614898 290382 615454
rect 289826 578898 290382 579454
rect 289826 542898 290382 543454
rect 289826 506898 290382 507454
rect 289826 470898 290382 471454
rect 289826 434898 290382 435454
rect 289826 398898 290382 399454
rect 293546 690618 294102 691174
rect 293546 654618 294102 655174
rect 293546 618618 294102 619174
rect 293546 582618 294102 583174
rect 293546 546618 294102 547174
rect 293546 510618 294102 511174
rect 293546 474618 294102 475174
rect 293546 438618 294102 439174
rect 293546 402618 294102 403174
rect 297266 694338 297822 694894
rect 297266 658338 297822 658894
rect 297266 622338 297822 622894
rect 297266 586338 297822 586894
rect 297266 550338 297822 550894
rect 297266 514338 297822 514894
rect 297266 478338 297822 478894
rect 297266 442338 297822 442894
rect 297266 406338 297822 406894
rect 228986 374058 229542 374614
rect 228986 338058 229542 338614
rect 228986 302058 229542 302614
rect 228986 266058 229542 266614
rect 228986 230058 229542 230614
rect 228986 194058 229542 194614
rect 228986 158058 229542 158614
rect 228986 122058 229542 122614
rect 228986 86058 229542 86614
rect 228986 50058 229542 50614
rect 228986 14058 229542 14614
rect 210986 -7622 211542 -7066
rect 235826 308898 236382 309454
rect 235826 272898 236382 273454
rect 235826 236898 236382 237454
rect 235826 200898 236382 201454
rect 235826 164898 236382 165454
rect 235826 128898 236382 129454
rect 235826 92898 236382 93454
rect 235826 56898 236382 57454
rect 235826 20898 236382 21454
rect 239250 363218 239486 363454
rect 239250 362898 239486 363134
rect 239546 312618 240102 313174
rect 239546 276618 240102 277174
rect 239546 240618 240102 241174
rect 239546 204618 240102 205174
rect 239546 168618 240102 169174
rect 243266 316338 243822 316894
rect 243266 280338 243822 280894
rect 243266 244338 243822 244894
rect 269970 363218 270206 363454
rect 269970 362898 270206 363134
rect 254610 345218 254846 345454
rect 254610 344898 254846 345134
rect 285330 345218 285566 345454
rect 285330 344898 285566 345134
rect 246986 320058 247542 320614
rect 246986 284058 247542 284614
rect 246986 248058 247542 248614
rect 243266 208338 243822 208894
rect 243266 172338 243822 172894
rect 239546 132618 240102 133174
rect 239546 96618 240102 97174
rect 239546 60618 240102 61174
rect 239546 24618 240102 25174
rect 235826 -1862 236382 -1306
rect 239546 -3782 240102 -3226
rect 243266 136338 243822 136894
rect 243266 100338 243822 100894
rect 243266 64338 243822 64894
rect 243266 28338 243822 28894
rect 243266 -5702 243822 -5146
rect 246986 212058 247542 212614
rect 246986 176058 247542 176614
rect 246986 140058 247542 140614
rect 246986 104058 247542 104614
rect 246986 68058 247542 68614
rect 246986 32058 247542 32614
rect 228986 -6662 229542 -6106
rect 253826 326898 254382 327454
rect 253826 290898 254382 291454
rect 253826 254898 254382 255454
rect 253826 218898 254382 219454
rect 253826 182898 254382 183454
rect 253826 146898 254382 147454
rect 253826 110898 254382 111454
rect 253826 74898 254382 75454
rect 253826 38898 254382 39454
rect 253826 2898 254382 3454
rect 253826 -902 254382 -346
rect 257546 330618 258102 331174
rect 257546 294618 258102 295174
rect 257546 258618 258102 259174
rect 257546 222618 258102 223174
rect 257546 186618 258102 187174
rect 257546 150618 258102 151174
rect 257546 114618 258102 115174
rect 257546 78618 258102 79174
rect 257546 42618 258102 43174
rect 257546 6618 258102 7174
rect 257546 -2822 258102 -2266
rect 261266 334338 261822 334894
rect 261266 298338 261822 298894
rect 261266 262338 261822 262894
rect 261266 226338 261822 226894
rect 261266 190338 261822 190894
rect 261266 154338 261822 154894
rect 261266 118338 261822 118894
rect 261266 82338 261822 82894
rect 261266 46338 261822 46894
rect 261266 10338 261822 10894
rect 261266 -4742 261822 -4186
rect 264986 302058 265542 302614
rect 264986 266058 265542 266614
rect 264986 230058 265542 230614
rect 264986 194058 265542 194614
rect 264986 158058 265542 158614
rect 264986 122058 265542 122614
rect 264986 86058 265542 86614
rect 264986 50058 265542 50614
rect 264986 14058 265542 14614
rect 246986 -7622 247542 -7066
rect 271826 308898 272382 309454
rect 271826 272898 272382 273454
rect 271826 236898 272382 237454
rect 271826 200898 272382 201454
rect 271826 164898 272382 165454
rect 271826 128898 272382 129454
rect 271826 92898 272382 93454
rect 271826 56898 272382 57454
rect 271826 20898 272382 21454
rect 271826 -1862 272382 -1306
rect 275546 312618 276102 313174
rect 275546 276618 276102 277174
rect 275546 240618 276102 241174
rect 275546 204618 276102 205174
rect 275546 168618 276102 169174
rect 275546 132618 276102 133174
rect 275546 96618 276102 97174
rect 275546 60618 276102 61174
rect 275546 24618 276102 25174
rect 275546 -3782 276102 -3226
rect 279266 316338 279822 316894
rect 279266 280338 279822 280894
rect 279266 244338 279822 244894
rect 279266 208338 279822 208894
rect 279266 172338 279822 172894
rect 279266 136338 279822 136894
rect 279266 100338 279822 100894
rect 279266 64338 279822 64894
rect 279266 28338 279822 28894
rect 279266 -5702 279822 -5146
rect 282986 320058 283542 320614
rect 282986 284058 283542 284614
rect 282986 248058 283542 248614
rect 282986 212058 283542 212614
rect 282986 176058 283542 176614
rect 282986 140058 283542 140614
rect 289826 326898 290382 327454
rect 289826 290898 290382 291454
rect 289826 254898 290382 255454
rect 289826 218898 290382 219454
rect 289826 182898 290382 183454
rect 289826 146898 290382 147454
rect 282986 104058 283542 104614
rect 282986 68058 283542 68614
rect 282986 32058 283542 32614
rect 264986 -6662 265542 -6106
rect 289826 110898 290382 111454
rect 289826 74898 290382 75454
rect 297266 370338 297822 370894
rect 293546 330618 294102 331174
rect 293546 294618 294102 295174
rect 293546 258618 294102 259174
rect 293546 222618 294102 223174
rect 293546 186618 294102 187174
rect 293546 150618 294102 151174
rect 293546 114618 294102 115174
rect 293546 78618 294102 79174
rect 289826 38898 290382 39454
rect 289826 2898 290382 3454
rect 289826 -902 290382 -346
rect 293546 42618 294102 43174
rect 293546 6618 294102 7174
rect 293546 -2822 294102 -2266
rect 297266 334338 297822 334894
rect 297266 298338 297822 298894
rect 297266 262338 297822 262894
rect 297266 226338 297822 226894
rect 297266 190338 297822 190894
rect 297266 154338 297822 154894
rect 297266 118338 297822 118894
rect 297266 82338 297822 82894
rect 297266 46338 297822 46894
rect 297266 10338 297822 10894
rect 297266 -4742 297822 -4186
rect 318986 711002 319542 711558
rect 315266 709082 315822 709638
rect 311546 707162 312102 707718
rect 300986 698058 301542 698614
rect 300986 662058 301542 662614
rect 300986 626058 301542 626614
rect 300986 590058 301542 590614
rect 300986 554058 301542 554614
rect 300986 518058 301542 518614
rect 300986 482058 301542 482614
rect 300986 446058 301542 446614
rect 300986 410058 301542 410614
rect 300986 374058 301542 374614
rect 300986 338058 301542 338614
rect 300986 302058 301542 302614
rect 300986 266058 301542 266614
rect 300986 230058 301542 230614
rect 300986 194058 301542 194614
rect 300986 158058 301542 158614
rect 300986 122058 301542 122614
rect 300986 86058 301542 86614
rect 300986 50058 301542 50614
rect 300986 14058 301542 14614
rect 282986 -7622 283542 -7066
rect 307826 705242 308382 705798
rect 307826 668898 308382 669454
rect 307826 632898 308382 633454
rect 307826 596898 308382 597454
rect 307826 560898 308382 561454
rect 307826 524898 308382 525454
rect 307826 488898 308382 489454
rect 307826 452898 308382 453454
rect 307826 416898 308382 417454
rect 307826 380898 308382 381454
rect 307826 344898 308382 345454
rect 307826 308898 308382 309454
rect 307826 272898 308382 273454
rect 307826 236898 308382 237454
rect 307826 200898 308382 201454
rect 307826 164898 308382 165454
rect 307826 128898 308382 129454
rect 307826 92898 308382 93454
rect 307826 56898 308382 57454
rect 307826 20898 308382 21454
rect 307826 -1862 308382 -1306
rect 311546 672618 312102 673174
rect 311546 636618 312102 637174
rect 311546 600618 312102 601174
rect 311546 564618 312102 565174
rect 311546 528618 312102 529174
rect 311546 492618 312102 493174
rect 311546 456618 312102 457174
rect 311546 420618 312102 421174
rect 311546 384618 312102 385174
rect 311546 348618 312102 349174
rect 311546 312618 312102 313174
rect 311546 276618 312102 277174
rect 311546 240618 312102 241174
rect 311546 204618 312102 205174
rect 311546 168618 312102 169174
rect 311546 132618 312102 133174
rect 311546 96618 312102 97174
rect 311546 60618 312102 61174
rect 311546 24618 312102 25174
rect 311546 -3782 312102 -3226
rect 315266 676338 315822 676894
rect 315266 640338 315822 640894
rect 315266 604338 315822 604894
rect 315266 568338 315822 568894
rect 315266 532338 315822 532894
rect 315266 496338 315822 496894
rect 315266 460338 315822 460894
rect 315266 424338 315822 424894
rect 315266 388338 315822 388894
rect 315266 352338 315822 352894
rect 315266 316338 315822 316894
rect 315266 280338 315822 280894
rect 315266 244338 315822 244894
rect 315266 208338 315822 208894
rect 315266 172338 315822 172894
rect 315266 136338 315822 136894
rect 315266 100338 315822 100894
rect 315266 64338 315822 64894
rect 315266 28338 315822 28894
rect 315266 -5702 315822 -5146
rect 336986 710042 337542 710598
rect 333266 708122 333822 708678
rect 329546 706202 330102 706758
rect 318986 680058 319542 680614
rect 318986 644058 319542 644614
rect 318986 608058 319542 608614
rect 318986 572058 319542 572614
rect 318986 536058 319542 536614
rect 318986 500058 319542 500614
rect 318986 464058 319542 464614
rect 318986 428058 319542 428614
rect 318986 392058 319542 392614
rect 318986 356058 319542 356614
rect 318986 320058 319542 320614
rect 318986 284058 319542 284614
rect 318986 248058 319542 248614
rect 318986 212058 319542 212614
rect 318986 176058 319542 176614
rect 318986 140058 319542 140614
rect 318986 104058 319542 104614
rect 318986 68058 319542 68614
rect 318986 32058 319542 32614
rect 300986 -6662 301542 -6106
rect 325826 704282 326382 704838
rect 325826 686898 326382 687454
rect 325826 650898 326382 651454
rect 325826 614898 326382 615454
rect 325826 578898 326382 579454
rect 325826 542898 326382 543454
rect 325826 506898 326382 507454
rect 325826 470898 326382 471454
rect 325826 434898 326382 435454
rect 325826 398898 326382 399454
rect 325826 362898 326382 363454
rect 325826 326898 326382 327454
rect 325826 290898 326382 291454
rect 325826 254898 326382 255454
rect 325826 218898 326382 219454
rect 325826 182898 326382 183454
rect 325826 146898 326382 147454
rect 325826 110898 326382 111454
rect 325826 74898 326382 75454
rect 325826 38898 326382 39454
rect 325826 2898 326382 3454
rect 325826 -902 326382 -346
rect 329546 690618 330102 691174
rect 329546 654618 330102 655174
rect 329546 618618 330102 619174
rect 329546 582618 330102 583174
rect 329546 546618 330102 547174
rect 329546 510618 330102 511174
rect 329546 474618 330102 475174
rect 329546 438618 330102 439174
rect 329546 402618 330102 403174
rect 329546 366618 330102 367174
rect 329546 330618 330102 331174
rect 329546 294618 330102 295174
rect 329546 258618 330102 259174
rect 329546 222618 330102 223174
rect 329546 186618 330102 187174
rect 329546 150618 330102 151174
rect 329546 114618 330102 115174
rect 329546 78618 330102 79174
rect 329546 42618 330102 43174
rect 329546 6618 330102 7174
rect 329546 -2822 330102 -2266
rect 333266 694338 333822 694894
rect 333266 658338 333822 658894
rect 333266 622338 333822 622894
rect 333266 586338 333822 586894
rect 333266 550338 333822 550894
rect 333266 514338 333822 514894
rect 333266 478338 333822 478894
rect 333266 442338 333822 442894
rect 333266 406338 333822 406894
rect 333266 370338 333822 370894
rect 333266 334338 333822 334894
rect 333266 298338 333822 298894
rect 333266 262338 333822 262894
rect 333266 226338 333822 226894
rect 333266 190338 333822 190894
rect 333266 154338 333822 154894
rect 333266 118338 333822 118894
rect 333266 82338 333822 82894
rect 333266 46338 333822 46894
rect 333266 10338 333822 10894
rect 333266 -4742 333822 -4186
rect 354986 711002 355542 711558
rect 351266 709082 351822 709638
rect 347546 707162 348102 707718
rect 336986 698058 337542 698614
rect 336986 662058 337542 662614
rect 336986 626058 337542 626614
rect 336986 590058 337542 590614
rect 336986 554058 337542 554614
rect 336986 518058 337542 518614
rect 336986 482058 337542 482614
rect 336986 446058 337542 446614
rect 336986 410058 337542 410614
rect 336986 374058 337542 374614
rect 336986 338058 337542 338614
rect 336986 302058 337542 302614
rect 336986 266058 337542 266614
rect 336986 230058 337542 230614
rect 336986 194058 337542 194614
rect 336986 158058 337542 158614
rect 336986 122058 337542 122614
rect 336986 86058 337542 86614
rect 336986 50058 337542 50614
rect 336986 14058 337542 14614
rect 318986 -7622 319542 -7066
rect 343826 705242 344382 705798
rect 343826 668898 344382 669454
rect 343826 632898 344382 633454
rect 343826 596898 344382 597454
rect 343826 560898 344382 561454
rect 343826 524898 344382 525454
rect 343826 488898 344382 489454
rect 343826 452898 344382 453454
rect 343826 416898 344382 417454
rect 343826 380898 344382 381454
rect 343826 344898 344382 345454
rect 343826 308898 344382 309454
rect 343826 272898 344382 273454
rect 343826 236898 344382 237454
rect 343826 200898 344382 201454
rect 343826 164898 344382 165454
rect 343826 128898 344382 129454
rect 343826 92898 344382 93454
rect 343826 56898 344382 57454
rect 343826 20898 344382 21454
rect 343826 -1862 344382 -1306
rect 347546 672618 348102 673174
rect 347546 636618 348102 637174
rect 347546 600618 348102 601174
rect 347546 564618 348102 565174
rect 347546 528618 348102 529174
rect 347546 492618 348102 493174
rect 347546 456618 348102 457174
rect 347546 420618 348102 421174
rect 347546 384618 348102 385174
rect 347546 348618 348102 349174
rect 347546 312618 348102 313174
rect 347546 276618 348102 277174
rect 347546 240618 348102 241174
rect 347546 204618 348102 205174
rect 347546 168618 348102 169174
rect 347546 132618 348102 133174
rect 347546 96618 348102 97174
rect 347546 60618 348102 61174
rect 347546 24618 348102 25174
rect 347546 -3782 348102 -3226
rect 351266 676338 351822 676894
rect 351266 640338 351822 640894
rect 351266 604338 351822 604894
rect 351266 568338 351822 568894
rect 351266 532338 351822 532894
rect 351266 496338 351822 496894
rect 351266 460338 351822 460894
rect 351266 424338 351822 424894
rect 351266 388338 351822 388894
rect 351266 352338 351822 352894
rect 351266 316338 351822 316894
rect 351266 280338 351822 280894
rect 351266 244338 351822 244894
rect 351266 208338 351822 208894
rect 351266 172338 351822 172894
rect 351266 136338 351822 136894
rect 351266 100338 351822 100894
rect 351266 64338 351822 64894
rect 351266 28338 351822 28894
rect 351266 -5702 351822 -5146
rect 372986 710042 373542 710598
rect 369266 708122 369822 708678
rect 365546 706202 366102 706758
rect 354986 680058 355542 680614
rect 354986 644058 355542 644614
rect 354986 608058 355542 608614
rect 354986 572058 355542 572614
rect 354986 536058 355542 536614
rect 354986 500058 355542 500614
rect 354986 464058 355542 464614
rect 354986 428058 355542 428614
rect 354986 392058 355542 392614
rect 354986 356058 355542 356614
rect 354986 320058 355542 320614
rect 354986 284058 355542 284614
rect 354986 248058 355542 248614
rect 354986 212058 355542 212614
rect 354986 176058 355542 176614
rect 354986 140058 355542 140614
rect 354986 104058 355542 104614
rect 354986 68058 355542 68614
rect 354986 32058 355542 32614
rect 336986 -6662 337542 -6106
rect 361826 704282 362382 704838
rect 361826 686898 362382 687454
rect 361826 650898 362382 651454
rect 361826 614898 362382 615454
rect 361826 578898 362382 579454
rect 361826 542898 362382 543454
rect 361826 506898 362382 507454
rect 361826 470898 362382 471454
rect 361826 434898 362382 435454
rect 361826 398898 362382 399454
rect 361826 362898 362382 363454
rect 361826 326898 362382 327454
rect 361826 290898 362382 291454
rect 361826 254898 362382 255454
rect 361826 218898 362382 219454
rect 361826 182898 362382 183454
rect 361826 146898 362382 147454
rect 361826 110898 362382 111454
rect 361826 74898 362382 75454
rect 361826 38898 362382 39454
rect 361826 2898 362382 3454
rect 361826 -902 362382 -346
rect 365546 690618 366102 691174
rect 365546 654618 366102 655174
rect 365546 618618 366102 619174
rect 365546 582618 366102 583174
rect 365546 546618 366102 547174
rect 365546 510618 366102 511174
rect 365546 474618 366102 475174
rect 365546 438618 366102 439174
rect 365546 402618 366102 403174
rect 365546 366618 366102 367174
rect 365546 330618 366102 331174
rect 365546 294618 366102 295174
rect 365546 258618 366102 259174
rect 365546 222618 366102 223174
rect 365546 186618 366102 187174
rect 365546 150618 366102 151174
rect 365546 114618 366102 115174
rect 365546 78618 366102 79174
rect 365546 42618 366102 43174
rect 365546 6618 366102 7174
rect 365546 -2822 366102 -2266
rect 369266 694338 369822 694894
rect 369266 658338 369822 658894
rect 369266 622338 369822 622894
rect 369266 586338 369822 586894
rect 369266 550338 369822 550894
rect 369266 514338 369822 514894
rect 369266 478338 369822 478894
rect 369266 442338 369822 442894
rect 369266 406338 369822 406894
rect 369266 370338 369822 370894
rect 369266 334338 369822 334894
rect 369266 298338 369822 298894
rect 369266 262338 369822 262894
rect 369266 226338 369822 226894
rect 369266 190338 369822 190894
rect 369266 154338 369822 154894
rect 369266 118338 369822 118894
rect 369266 82338 369822 82894
rect 369266 46338 369822 46894
rect 369266 10338 369822 10894
rect 369266 -4742 369822 -4186
rect 390986 711002 391542 711558
rect 387266 709082 387822 709638
rect 383546 707162 384102 707718
rect 372986 698058 373542 698614
rect 372986 662058 373542 662614
rect 372986 626058 373542 626614
rect 372986 590058 373542 590614
rect 372986 554058 373542 554614
rect 372986 518058 373542 518614
rect 372986 482058 373542 482614
rect 372986 446058 373542 446614
rect 372986 410058 373542 410614
rect 372986 374058 373542 374614
rect 372986 338058 373542 338614
rect 372986 302058 373542 302614
rect 372986 266058 373542 266614
rect 372986 230058 373542 230614
rect 372986 194058 373542 194614
rect 372986 158058 373542 158614
rect 372986 122058 373542 122614
rect 372986 86058 373542 86614
rect 372986 50058 373542 50614
rect 372986 14058 373542 14614
rect 354986 -7622 355542 -7066
rect 379826 705242 380382 705798
rect 379826 668898 380382 669454
rect 379826 632898 380382 633454
rect 379826 596898 380382 597454
rect 379826 560898 380382 561454
rect 379826 524898 380382 525454
rect 379826 488898 380382 489454
rect 379826 452898 380382 453454
rect 379826 416898 380382 417454
rect 379826 380898 380382 381454
rect 379826 344898 380382 345454
rect 379826 308898 380382 309454
rect 379826 272898 380382 273454
rect 379826 236898 380382 237454
rect 379826 200898 380382 201454
rect 379826 164898 380382 165454
rect 379826 128898 380382 129454
rect 379826 92898 380382 93454
rect 379826 56898 380382 57454
rect 379826 20898 380382 21454
rect 379826 -1862 380382 -1306
rect 383546 672618 384102 673174
rect 383546 636618 384102 637174
rect 383546 600618 384102 601174
rect 383546 564618 384102 565174
rect 383546 528618 384102 529174
rect 383546 492618 384102 493174
rect 383546 456618 384102 457174
rect 383546 420618 384102 421174
rect 383546 384618 384102 385174
rect 383546 348618 384102 349174
rect 383546 312618 384102 313174
rect 383546 276618 384102 277174
rect 383546 240618 384102 241174
rect 383546 204618 384102 205174
rect 383546 168618 384102 169174
rect 383546 132618 384102 133174
rect 383546 96618 384102 97174
rect 383546 60618 384102 61174
rect 383546 24618 384102 25174
rect 383546 -3782 384102 -3226
rect 387266 676338 387822 676894
rect 387266 640338 387822 640894
rect 387266 604338 387822 604894
rect 387266 568338 387822 568894
rect 387266 532338 387822 532894
rect 387266 496338 387822 496894
rect 387266 460338 387822 460894
rect 387266 424338 387822 424894
rect 387266 388338 387822 388894
rect 387266 352338 387822 352894
rect 387266 316338 387822 316894
rect 387266 280338 387822 280894
rect 387266 244338 387822 244894
rect 387266 208338 387822 208894
rect 387266 172338 387822 172894
rect 387266 136338 387822 136894
rect 387266 100338 387822 100894
rect 387266 64338 387822 64894
rect 387266 28338 387822 28894
rect 387266 -5702 387822 -5146
rect 408986 710042 409542 710598
rect 405266 708122 405822 708678
rect 401546 706202 402102 706758
rect 390986 680058 391542 680614
rect 390986 644058 391542 644614
rect 390986 608058 391542 608614
rect 390986 572058 391542 572614
rect 390986 536058 391542 536614
rect 390986 500058 391542 500614
rect 390986 464058 391542 464614
rect 390986 428058 391542 428614
rect 390986 392058 391542 392614
rect 390986 356058 391542 356614
rect 390986 320058 391542 320614
rect 390986 284058 391542 284614
rect 390986 248058 391542 248614
rect 390986 212058 391542 212614
rect 390986 176058 391542 176614
rect 390986 140058 391542 140614
rect 390986 104058 391542 104614
rect 390986 68058 391542 68614
rect 390986 32058 391542 32614
rect 372986 -6662 373542 -6106
rect 397826 704282 398382 704838
rect 397826 686898 398382 687454
rect 397826 650898 398382 651454
rect 397826 614898 398382 615454
rect 397826 578898 398382 579454
rect 397826 542898 398382 543454
rect 397826 506898 398382 507454
rect 397826 470898 398382 471454
rect 397826 434898 398382 435454
rect 397826 398898 398382 399454
rect 397826 362898 398382 363454
rect 397826 326898 398382 327454
rect 397826 290898 398382 291454
rect 397826 254898 398382 255454
rect 397826 218898 398382 219454
rect 397826 182898 398382 183454
rect 397826 146898 398382 147454
rect 397826 110898 398382 111454
rect 397826 74898 398382 75454
rect 397826 38898 398382 39454
rect 397826 2898 398382 3454
rect 397826 -902 398382 -346
rect 401546 690618 402102 691174
rect 401546 654618 402102 655174
rect 401546 618618 402102 619174
rect 401546 582618 402102 583174
rect 401546 546618 402102 547174
rect 401546 510618 402102 511174
rect 401546 474618 402102 475174
rect 401546 438618 402102 439174
rect 401546 402618 402102 403174
rect 401546 366618 402102 367174
rect 401546 330618 402102 331174
rect 401546 294618 402102 295174
rect 401546 258618 402102 259174
rect 401546 222618 402102 223174
rect 401546 186618 402102 187174
rect 401546 150618 402102 151174
rect 401546 114618 402102 115174
rect 401546 78618 402102 79174
rect 401546 42618 402102 43174
rect 401546 6618 402102 7174
rect 401546 -2822 402102 -2266
rect 405266 694338 405822 694894
rect 405266 658338 405822 658894
rect 405266 622338 405822 622894
rect 405266 586338 405822 586894
rect 405266 550338 405822 550894
rect 405266 514338 405822 514894
rect 405266 478338 405822 478894
rect 405266 442338 405822 442894
rect 405266 406338 405822 406894
rect 405266 370338 405822 370894
rect 405266 334338 405822 334894
rect 405266 298338 405822 298894
rect 405266 262338 405822 262894
rect 405266 226338 405822 226894
rect 405266 190338 405822 190894
rect 405266 154338 405822 154894
rect 405266 118338 405822 118894
rect 405266 82338 405822 82894
rect 405266 46338 405822 46894
rect 405266 10338 405822 10894
rect 405266 -4742 405822 -4186
rect 426986 711002 427542 711558
rect 423266 709082 423822 709638
rect 419546 707162 420102 707718
rect 408986 698058 409542 698614
rect 408986 662058 409542 662614
rect 408986 626058 409542 626614
rect 408986 590058 409542 590614
rect 408986 554058 409542 554614
rect 408986 518058 409542 518614
rect 408986 482058 409542 482614
rect 408986 446058 409542 446614
rect 408986 410058 409542 410614
rect 408986 374058 409542 374614
rect 408986 338058 409542 338614
rect 408986 302058 409542 302614
rect 408986 266058 409542 266614
rect 408986 230058 409542 230614
rect 408986 194058 409542 194614
rect 408986 158058 409542 158614
rect 408986 122058 409542 122614
rect 408986 86058 409542 86614
rect 408986 50058 409542 50614
rect 408986 14058 409542 14614
rect 390986 -7622 391542 -7066
rect 415826 705242 416382 705798
rect 415826 668898 416382 669454
rect 415826 632898 416382 633454
rect 415826 596898 416382 597454
rect 415826 560898 416382 561454
rect 415826 524898 416382 525454
rect 415826 488898 416382 489454
rect 415826 452898 416382 453454
rect 415826 416898 416382 417454
rect 415826 380898 416382 381454
rect 415826 344898 416382 345454
rect 415826 308898 416382 309454
rect 415826 272898 416382 273454
rect 415826 236898 416382 237454
rect 415826 200898 416382 201454
rect 415826 164898 416382 165454
rect 415826 128898 416382 129454
rect 415826 92898 416382 93454
rect 415826 56898 416382 57454
rect 415826 20898 416382 21454
rect 415826 -1862 416382 -1306
rect 419546 672618 420102 673174
rect 419546 636618 420102 637174
rect 419546 600618 420102 601174
rect 419546 564618 420102 565174
rect 419546 528618 420102 529174
rect 419546 492618 420102 493174
rect 419546 456618 420102 457174
rect 419546 420618 420102 421174
rect 419546 384618 420102 385174
rect 419546 348618 420102 349174
rect 419546 312618 420102 313174
rect 419546 276618 420102 277174
rect 419546 240618 420102 241174
rect 419546 204618 420102 205174
rect 419546 168618 420102 169174
rect 419546 132618 420102 133174
rect 419546 96618 420102 97174
rect 419546 60618 420102 61174
rect 419546 24618 420102 25174
rect 419546 -3782 420102 -3226
rect 423266 676338 423822 676894
rect 423266 640338 423822 640894
rect 423266 604338 423822 604894
rect 423266 568338 423822 568894
rect 423266 532338 423822 532894
rect 423266 496338 423822 496894
rect 423266 460338 423822 460894
rect 423266 424338 423822 424894
rect 423266 388338 423822 388894
rect 423266 352338 423822 352894
rect 423266 316338 423822 316894
rect 423266 280338 423822 280894
rect 423266 244338 423822 244894
rect 423266 208338 423822 208894
rect 423266 172338 423822 172894
rect 423266 136338 423822 136894
rect 423266 100338 423822 100894
rect 423266 64338 423822 64894
rect 423266 28338 423822 28894
rect 423266 -5702 423822 -5146
rect 444986 710042 445542 710598
rect 441266 708122 441822 708678
rect 437546 706202 438102 706758
rect 426986 680058 427542 680614
rect 426986 644058 427542 644614
rect 426986 608058 427542 608614
rect 426986 572058 427542 572614
rect 426986 536058 427542 536614
rect 426986 500058 427542 500614
rect 426986 464058 427542 464614
rect 426986 428058 427542 428614
rect 426986 392058 427542 392614
rect 426986 356058 427542 356614
rect 426986 320058 427542 320614
rect 426986 284058 427542 284614
rect 426986 248058 427542 248614
rect 426986 212058 427542 212614
rect 426986 176058 427542 176614
rect 426986 140058 427542 140614
rect 426986 104058 427542 104614
rect 426986 68058 427542 68614
rect 426986 32058 427542 32614
rect 408986 -6662 409542 -6106
rect 433826 704282 434382 704838
rect 433826 686898 434382 687454
rect 433826 650898 434382 651454
rect 433826 614898 434382 615454
rect 433826 578898 434382 579454
rect 433826 542898 434382 543454
rect 433826 506898 434382 507454
rect 433826 470898 434382 471454
rect 433826 434898 434382 435454
rect 433826 398898 434382 399454
rect 433826 362898 434382 363454
rect 433826 326898 434382 327454
rect 433826 290898 434382 291454
rect 433826 254898 434382 255454
rect 433826 218898 434382 219454
rect 433826 182898 434382 183454
rect 433826 146898 434382 147454
rect 433826 110898 434382 111454
rect 433826 74898 434382 75454
rect 433826 38898 434382 39454
rect 433826 2898 434382 3454
rect 433826 -902 434382 -346
rect 437546 690618 438102 691174
rect 437546 654618 438102 655174
rect 437546 618618 438102 619174
rect 437546 582618 438102 583174
rect 437546 546618 438102 547174
rect 437546 510618 438102 511174
rect 437546 474618 438102 475174
rect 437546 438618 438102 439174
rect 437546 402618 438102 403174
rect 437546 366618 438102 367174
rect 437546 330618 438102 331174
rect 437546 294618 438102 295174
rect 437546 258618 438102 259174
rect 437546 222618 438102 223174
rect 437546 186618 438102 187174
rect 437546 150618 438102 151174
rect 437546 114618 438102 115174
rect 437546 78618 438102 79174
rect 437546 42618 438102 43174
rect 437546 6618 438102 7174
rect 437546 -2822 438102 -2266
rect 441266 694338 441822 694894
rect 441266 658338 441822 658894
rect 441266 622338 441822 622894
rect 441266 586338 441822 586894
rect 441266 550338 441822 550894
rect 441266 514338 441822 514894
rect 441266 478338 441822 478894
rect 441266 442338 441822 442894
rect 441266 406338 441822 406894
rect 441266 370338 441822 370894
rect 441266 334338 441822 334894
rect 441266 298338 441822 298894
rect 441266 262338 441822 262894
rect 441266 226338 441822 226894
rect 441266 190338 441822 190894
rect 441266 154338 441822 154894
rect 441266 118338 441822 118894
rect 441266 82338 441822 82894
rect 441266 46338 441822 46894
rect 441266 10338 441822 10894
rect 441266 -4742 441822 -4186
rect 462986 711002 463542 711558
rect 459266 709082 459822 709638
rect 455546 707162 456102 707718
rect 444986 698058 445542 698614
rect 444986 662058 445542 662614
rect 444986 626058 445542 626614
rect 444986 590058 445542 590614
rect 444986 554058 445542 554614
rect 444986 518058 445542 518614
rect 444986 482058 445542 482614
rect 444986 446058 445542 446614
rect 444986 410058 445542 410614
rect 444986 374058 445542 374614
rect 444986 338058 445542 338614
rect 444986 302058 445542 302614
rect 444986 266058 445542 266614
rect 444986 230058 445542 230614
rect 444986 194058 445542 194614
rect 444986 158058 445542 158614
rect 444986 122058 445542 122614
rect 444986 86058 445542 86614
rect 444986 50058 445542 50614
rect 444986 14058 445542 14614
rect 426986 -7622 427542 -7066
rect 451826 705242 452382 705798
rect 451826 668898 452382 669454
rect 451826 632898 452382 633454
rect 451826 596898 452382 597454
rect 451826 560898 452382 561454
rect 451826 524898 452382 525454
rect 451826 488898 452382 489454
rect 451826 452898 452382 453454
rect 451826 416898 452382 417454
rect 451826 380898 452382 381454
rect 451826 344898 452382 345454
rect 451826 308898 452382 309454
rect 451826 272898 452382 273454
rect 451826 236898 452382 237454
rect 451826 200898 452382 201454
rect 451826 164898 452382 165454
rect 451826 128898 452382 129454
rect 451826 92898 452382 93454
rect 451826 56898 452382 57454
rect 451826 20898 452382 21454
rect 451826 -1862 452382 -1306
rect 455546 672618 456102 673174
rect 455546 636618 456102 637174
rect 455546 600618 456102 601174
rect 455546 564618 456102 565174
rect 455546 528618 456102 529174
rect 455546 492618 456102 493174
rect 455546 456618 456102 457174
rect 455546 420618 456102 421174
rect 455546 384618 456102 385174
rect 455546 348618 456102 349174
rect 455546 312618 456102 313174
rect 455546 276618 456102 277174
rect 455546 240618 456102 241174
rect 455546 204618 456102 205174
rect 455546 168618 456102 169174
rect 455546 132618 456102 133174
rect 455546 96618 456102 97174
rect 455546 60618 456102 61174
rect 455546 24618 456102 25174
rect 455546 -3782 456102 -3226
rect 459266 676338 459822 676894
rect 459266 640338 459822 640894
rect 459266 604338 459822 604894
rect 459266 568338 459822 568894
rect 459266 532338 459822 532894
rect 459266 496338 459822 496894
rect 459266 460338 459822 460894
rect 459266 424338 459822 424894
rect 459266 388338 459822 388894
rect 459266 352338 459822 352894
rect 459266 316338 459822 316894
rect 459266 280338 459822 280894
rect 459266 244338 459822 244894
rect 459266 208338 459822 208894
rect 459266 172338 459822 172894
rect 459266 136338 459822 136894
rect 459266 100338 459822 100894
rect 459266 64338 459822 64894
rect 459266 28338 459822 28894
rect 459266 -5702 459822 -5146
rect 480986 710042 481542 710598
rect 477266 708122 477822 708678
rect 473546 706202 474102 706758
rect 462986 680058 463542 680614
rect 462986 644058 463542 644614
rect 462986 608058 463542 608614
rect 462986 572058 463542 572614
rect 462986 536058 463542 536614
rect 462986 500058 463542 500614
rect 462986 464058 463542 464614
rect 462986 428058 463542 428614
rect 462986 392058 463542 392614
rect 462986 356058 463542 356614
rect 462986 320058 463542 320614
rect 462986 284058 463542 284614
rect 462986 248058 463542 248614
rect 462986 212058 463542 212614
rect 462986 176058 463542 176614
rect 462986 140058 463542 140614
rect 462986 104058 463542 104614
rect 462986 68058 463542 68614
rect 462986 32058 463542 32614
rect 444986 -6662 445542 -6106
rect 469826 704282 470382 704838
rect 469826 686898 470382 687454
rect 469826 650898 470382 651454
rect 469826 614898 470382 615454
rect 469826 578898 470382 579454
rect 469826 542898 470382 543454
rect 469826 506898 470382 507454
rect 469826 470898 470382 471454
rect 469826 434898 470382 435454
rect 469826 398898 470382 399454
rect 469826 362898 470382 363454
rect 469826 326898 470382 327454
rect 469826 290898 470382 291454
rect 469826 254898 470382 255454
rect 469826 218898 470382 219454
rect 469826 182898 470382 183454
rect 469826 146898 470382 147454
rect 469826 110898 470382 111454
rect 469826 74898 470382 75454
rect 469826 38898 470382 39454
rect 469826 2898 470382 3454
rect 469826 -902 470382 -346
rect 473546 690618 474102 691174
rect 473546 654618 474102 655174
rect 473546 618618 474102 619174
rect 473546 582618 474102 583174
rect 473546 546618 474102 547174
rect 473546 510618 474102 511174
rect 473546 474618 474102 475174
rect 473546 438618 474102 439174
rect 473546 402618 474102 403174
rect 473546 366618 474102 367174
rect 473546 330618 474102 331174
rect 473546 294618 474102 295174
rect 473546 258618 474102 259174
rect 473546 222618 474102 223174
rect 473546 186618 474102 187174
rect 473546 150618 474102 151174
rect 473546 114618 474102 115174
rect 473546 78618 474102 79174
rect 473546 42618 474102 43174
rect 473546 6618 474102 7174
rect 473546 -2822 474102 -2266
rect 477266 694338 477822 694894
rect 477266 658338 477822 658894
rect 477266 622338 477822 622894
rect 477266 586338 477822 586894
rect 477266 550338 477822 550894
rect 477266 514338 477822 514894
rect 477266 478338 477822 478894
rect 477266 442338 477822 442894
rect 477266 406338 477822 406894
rect 477266 370338 477822 370894
rect 477266 334338 477822 334894
rect 477266 298338 477822 298894
rect 477266 262338 477822 262894
rect 477266 226338 477822 226894
rect 477266 190338 477822 190894
rect 477266 154338 477822 154894
rect 477266 118338 477822 118894
rect 477266 82338 477822 82894
rect 477266 46338 477822 46894
rect 477266 10338 477822 10894
rect 477266 -4742 477822 -4186
rect 498986 711002 499542 711558
rect 495266 709082 495822 709638
rect 491546 707162 492102 707718
rect 480986 698058 481542 698614
rect 480986 662058 481542 662614
rect 480986 626058 481542 626614
rect 480986 590058 481542 590614
rect 480986 554058 481542 554614
rect 480986 518058 481542 518614
rect 480986 482058 481542 482614
rect 480986 446058 481542 446614
rect 480986 410058 481542 410614
rect 480986 374058 481542 374614
rect 480986 338058 481542 338614
rect 480986 302058 481542 302614
rect 480986 266058 481542 266614
rect 480986 230058 481542 230614
rect 480986 194058 481542 194614
rect 480986 158058 481542 158614
rect 480986 122058 481542 122614
rect 480986 86058 481542 86614
rect 480986 50058 481542 50614
rect 480986 14058 481542 14614
rect 462986 -7622 463542 -7066
rect 487826 705242 488382 705798
rect 487826 668898 488382 669454
rect 487826 632898 488382 633454
rect 487826 596898 488382 597454
rect 487826 560898 488382 561454
rect 487826 524898 488382 525454
rect 487826 488898 488382 489454
rect 487826 452898 488382 453454
rect 487826 416898 488382 417454
rect 487826 380898 488382 381454
rect 487826 344898 488382 345454
rect 487826 308898 488382 309454
rect 487826 272898 488382 273454
rect 487826 236898 488382 237454
rect 487826 200898 488382 201454
rect 487826 164898 488382 165454
rect 487826 128898 488382 129454
rect 487826 92898 488382 93454
rect 487826 56898 488382 57454
rect 487826 20898 488382 21454
rect 487826 -1862 488382 -1306
rect 491546 672618 492102 673174
rect 491546 636618 492102 637174
rect 491546 600618 492102 601174
rect 491546 564618 492102 565174
rect 491546 528618 492102 529174
rect 491546 492618 492102 493174
rect 491546 456618 492102 457174
rect 491546 420618 492102 421174
rect 491546 384618 492102 385174
rect 491546 348618 492102 349174
rect 491546 312618 492102 313174
rect 491546 276618 492102 277174
rect 491546 240618 492102 241174
rect 491546 204618 492102 205174
rect 491546 168618 492102 169174
rect 491546 132618 492102 133174
rect 491546 96618 492102 97174
rect 491546 60618 492102 61174
rect 491546 24618 492102 25174
rect 491546 -3782 492102 -3226
rect 495266 676338 495822 676894
rect 495266 640338 495822 640894
rect 495266 604338 495822 604894
rect 495266 568338 495822 568894
rect 495266 532338 495822 532894
rect 495266 496338 495822 496894
rect 495266 460338 495822 460894
rect 495266 424338 495822 424894
rect 495266 388338 495822 388894
rect 495266 352338 495822 352894
rect 495266 316338 495822 316894
rect 495266 280338 495822 280894
rect 495266 244338 495822 244894
rect 495266 208338 495822 208894
rect 495266 172338 495822 172894
rect 495266 136338 495822 136894
rect 495266 100338 495822 100894
rect 495266 64338 495822 64894
rect 495266 28338 495822 28894
rect 495266 -5702 495822 -5146
rect 516986 710042 517542 710598
rect 513266 708122 513822 708678
rect 509546 706202 510102 706758
rect 498986 680058 499542 680614
rect 498986 644058 499542 644614
rect 498986 608058 499542 608614
rect 498986 572058 499542 572614
rect 498986 536058 499542 536614
rect 498986 500058 499542 500614
rect 498986 464058 499542 464614
rect 498986 428058 499542 428614
rect 498986 392058 499542 392614
rect 498986 356058 499542 356614
rect 498986 320058 499542 320614
rect 498986 284058 499542 284614
rect 498986 248058 499542 248614
rect 498986 212058 499542 212614
rect 498986 176058 499542 176614
rect 498986 140058 499542 140614
rect 498986 104058 499542 104614
rect 498986 68058 499542 68614
rect 498986 32058 499542 32614
rect 480986 -6662 481542 -6106
rect 505826 704282 506382 704838
rect 505826 686898 506382 687454
rect 505826 650898 506382 651454
rect 505826 614898 506382 615454
rect 505826 578898 506382 579454
rect 505826 542898 506382 543454
rect 505826 506898 506382 507454
rect 505826 470898 506382 471454
rect 505826 434898 506382 435454
rect 505826 398898 506382 399454
rect 505826 362898 506382 363454
rect 505826 326898 506382 327454
rect 505826 290898 506382 291454
rect 505826 254898 506382 255454
rect 505826 218898 506382 219454
rect 505826 182898 506382 183454
rect 505826 146898 506382 147454
rect 505826 110898 506382 111454
rect 505826 74898 506382 75454
rect 505826 38898 506382 39454
rect 505826 2898 506382 3454
rect 505826 -902 506382 -346
rect 509546 690618 510102 691174
rect 509546 654618 510102 655174
rect 509546 618618 510102 619174
rect 509546 582618 510102 583174
rect 509546 546618 510102 547174
rect 509546 510618 510102 511174
rect 509546 474618 510102 475174
rect 509546 438618 510102 439174
rect 509546 402618 510102 403174
rect 509546 366618 510102 367174
rect 509546 330618 510102 331174
rect 509546 294618 510102 295174
rect 509546 258618 510102 259174
rect 509546 222618 510102 223174
rect 509546 186618 510102 187174
rect 509546 150618 510102 151174
rect 509546 114618 510102 115174
rect 509546 78618 510102 79174
rect 509546 42618 510102 43174
rect 509546 6618 510102 7174
rect 509546 -2822 510102 -2266
rect 513266 694338 513822 694894
rect 513266 658338 513822 658894
rect 513266 622338 513822 622894
rect 513266 586338 513822 586894
rect 513266 550338 513822 550894
rect 513266 514338 513822 514894
rect 513266 478338 513822 478894
rect 513266 442338 513822 442894
rect 513266 406338 513822 406894
rect 513266 370338 513822 370894
rect 513266 334338 513822 334894
rect 513266 298338 513822 298894
rect 513266 262338 513822 262894
rect 513266 226338 513822 226894
rect 513266 190338 513822 190894
rect 513266 154338 513822 154894
rect 513266 118338 513822 118894
rect 513266 82338 513822 82894
rect 513266 46338 513822 46894
rect 513266 10338 513822 10894
rect 513266 -4742 513822 -4186
rect 534986 711002 535542 711558
rect 531266 709082 531822 709638
rect 527546 707162 528102 707718
rect 516986 698058 517542 698614
rect 516986 662058 517542 662614
rect 516986 626058 517542 626614
rect 516986 590058 517542 590614
rect 516986 554058 517542 554614
rect 516986 518058 517542 518614
rect 516986 482058 517542 482614
rect 516986 446058 517542 446614
rect 516986 410058 517542 410614
rect 516986 374058 517542 374614
rect 516986 338058 517542 338614
rect 516986 302058 517542 302614
rect 516986 266058 517542 266614
rect 516986 230058 517542 230614
rect 516986 194058 517542 194614
rect 516986 158058 517542 158614
rect 516986 122058 517542 122614
rect 516986 86058 517542 86614
rect 516986 50058 517542 50614
rect 516986 14058 517542 14614
rect 498986 -7622 499542 -7066
rect 523826 705242 524382 705798
rect 523826 668898 524382 669454
rect 523826 632898 524382 633454
rect 523826 596898 524382 597454
rect 523826 560898 524382 561454
rect 523826 524898 524382 525454
rect 523826 488898 524382 489454
rect 523826 452898 524382 453454
rect 523826 416898 524382 417454
rect 523826 380898 524382 381454
rect 523826 344898 524382 345454
rect 523826 308898 524382 309454
rect 523826 272898 524382 273454
rect 523826 236898 524382 237454
rect 523826 200898 524382 201454
rect 523826 164898 524382 165454
rect 523826 128898 524382 129454
rect 523826 92898 524382 93454
rect 523826 56898 524382 57454
rect 523826 20898 524382 21454
rect 523826 -1862 524382 -1306
rect 527546 672618 528102 673174
rect 527546 636618 528102 637174
rect 527546 600618 528102 601174
rect 527546 564618 528102 565174
rect 527546 528618 528102 529174
rect 527546 492618 528102 493174
rect 527546 456618 528102 457174
rect 527546 420618 528102 421174
rect 527546 384618 528102 385174
rect 527546 348618 528102 349174
rect 527546 312618 528102 313174
rect 527546 276618 528102 277174
rect 527546 240618 528102 241174
rect 527546 204618 528102 205174
rect 527546 168618 528102 169174
rect 527546 132618 528102 133174
rect 527546 96618 528102 97174
rect 527546 60618 528102 61174
rect 527546 24618 528102 25174
rect 527546 -3782 528102 -3226
rect 531266 676338 531822 676894
rect 531266 640338 531822 640894
rect 531266 604338 531822 604894
rect 531266 568338 531822 568894
rect 531266 532338 531822 532894
rect 531266 496338 531822 496894
rect 531266 460338 531822 460894
rect 531266 424338 531822 424894
rect 531266 388338 531822 388894
rect 531266 352338 531822 352894
rect 531266 316338 531822 316894
rect 531266 280338 531822 280894
rect 531266 244338 531822 244894
rect 531266 208338 531822 208894
rect 531266 172338 531822 172894
rect 531266 136338 531822 136894
rect 531266 100338 531822 100894
rect 531266 64338 531822 64894
rect 531266 28338 531822 28894
rect 531266 -5702 531822 -5146
rect 552986 710042 553542 710598
rect 549266 708122 549822 708678
rect 545546 706202 546102 706758
rect 534986 680058 535542 680614
rect 534986 644058 535542 644614
rect 534986 608058 535542 608614
rect 534986 572058 535542 572614
rect 534986 536058 535542 536614
rect 534986 500058 535542 500614
rect 534986 464058 535542 464614
rect 534986 428058 535542 428614
rect 534986 392058 535542 392614
rect 534986 356058 535542 356614
rect 534986 320058 535542 320614
rect 534986 284058 535542 284614
rect 534986 248058 535542 248614
rect 534986 212058 535542 212614
rect 534986 176058 535542 176614
rect 534986 140058 535542 140614
rect 534986 104058 535542 104614
rect 534986 68058 535542 68614
rect 534986 32058 535542 32614
rect 516986 -6662 517542 -6106
rect 541826 704282 542382 704838
rect 541826 686898 542382 687454
rect 541826 650898 542382 651454
rect 541826 614898 542382 615454
rect 541826 578898 542382 579454
rect 541826 542898 542382 543454
rect 541826 506898 542382 507454
rect 541826 470898 542382 471454
rect 541826 434898 542382 435454
rect 541826 398898 542382 399454
rect 541826 362898 542382 363454
rect 541826 326898 542382 327454
rect 541826 290898 542382 291454
rect 541826 254898 542382 255454
rect 541826 218898 542382 219454
rect 541826 182898 542382 183454
rect 541826 146898 542382 147454
rect 541826 110898 542382 111454
rect 541826 74898 542382 75454
rect 541826 38898 542382 39454
rect 541826 2898 542382 3454
rect 541826 -902 542382 -346
rect 545546 690618 546102 691174
rect 545546 654618 546102 655174
rect 545546 618618 546102 619174
rect 545546 582618 546102 583174
rect 545546 546618 546102 547174
rect 545546 510618 546102 511174
rect 545546 474618 546102 475174
rect 545546 438618 546102 439174
rect 545546 402618 546102 403174
rect 545546 366618 546102 367174
rect 545546 330618 546102 331174
rect 545546 294618 546102 295174
rect 545546 258618 546102 259174
rect 545546 222618 546102 223174
rect 545546 186618 546102 187174
rect 545546 150618 546102 151174
rect 545546 114618 546102 115174
rect 545546 78618 546102 79174
rect 545546 42618 546102 43174
rect 545546 6618 546102 7174
rect 545546 -2822 546102 -2266
rect 549266 694338 549822 694894
rect 549266 658338 549822 658894
rect 549266 622338 549822 622894
rect 549266 586338 549822 586894
rect 549266 550338 549822 550894
rect 549266 514338 549822 514894
rect 549266 478338 549822 478894
rect 549266 442338 549822 442894
rect 549266 406338 549822 406894
rect 549266 370338 549822 370894
rect 549266 334338 549822 334894
rect 549266 298338 549822 298894
rect 549266 262338 549822 262894
rect 549266 226338 549822 226894
rect 549266 190338 549822 190894
rect 549266 154338 549822 154894
rect 549266 118338 549822 118894
rect 549266 82338 549822 82894
rect 549266 46338 549822 46894
rect 549266 10338 549822 10894
rect 549266 -4742 549822 -4186
rect 570986 711002 571542 711558
rect 567266 709082 567822 709638
rect 563546 707162 564102 707718
rect 552986 698058 553542 698614
rect 552986 662058 553542 662614
rect 552986 626058 553542 626614
rect 552986 590058 553542 590614
rect 552986 554058 553542 554614
rect 552986 518058 553542 518614
rect 552986 482058 553542 482614
rect 552986 446058 553542 446614
rect 552986 410058 553542 410614
rect 552986 374058 553542 374614
rect 552986 338058 553542 338614
rect 552986 302058 553542 302614
rect 552986 266058 553542 266614
rect 552986 230058 553542 230614
rect 552986 194058 553542 194614
rect 552986 158058 553542 158614
rect 552986 122058 553542 122614
rect 552986 86058 553542 86614
rect 552986 50058 553542 50614
rect 552986 14058 553542 14614
rect 534986 -7622 535542 -7066
rect 559826 705242 560382 705798
rect 559826 668898 560382 669454
rect 559826 632898 560382 633454
rect 559826 596898 560382 597454
rect 559826 560898 560382 561454
rect 559826 524898 560382 525454
rect 559826 488898 560382 489454
rect 559826 452898 560382 453454
rect 559826 416898 560382 417454
rect 559826 380898 560382 381454
rect 559826 344898 560382 345454
rect 559826 308898 560382 309454
rect 559826 272898 560382 273454
rect 559826 236898 560382 237454
rect 559826 200898 560382 201454
rect 559826 164898 560382 165454
rect 559826 128898 560382 129454
rect 559826 92898 560382 93454
rect 559826 56898 560382 57454
rect 559826 20898 560382 21454
rect 559826 -1862 560382 -1306
rect 563546 672618 564102 673174
rect 563546 636618 564102 637174
rect 563546 600618 564102 601174
rect 563546 564618 564102 565174
rect 563546 528618 564102 529174
rect 563546 492618 564102 493174
rect 563546 456618 564102 457174
rect 563546 420618 564102 421174
rect 563546 384618 564102 385174
rect 563546 348618 564102 349174
rect 563546 312618 564102 313174
rect 563546 276618 564102 277174
rect 563546 240618 564102 241174
rect 563546 204618 564102 205174
rect 563546 168618 564102 169174
rect 563546 132618 564102 133174
rect 563546 96618 564102 97174
rect 563546 60618 564102 61174
rect 563546 24618 564102 25174
rect 563546 -3782 564102 -3226
rect 567266 676338 567822 676894
rect 567266 640338 567822 640894
rect 567266 604338 567822 604894
rect 567266 568338 567822 568894
rect 567266 532338 567822 532894
rect 567266 496338 567822 496894
rect 567266 460338 567822 460894
rect 567266 424338 567822 424894
rect 567266 388338 567822 388894
rect 567266 352338 567822 352894
rect 567266 316338 567822 316894
rect 567266 280338 567822 280894
rect 567266 244338 567822 244894
rect 567266 208338 567822 208894
rect 567266 172338 567822 172894
rect 567266 136338 567822 136894
rect 567266 100338 567822 100894
rect 567266 64338 567822 64894
rect 567266 28338 567822 28894
rect 567266 -5702 567822 -5146
rect 592062 711002 592618 711558
rect 591102 710042 591658 710598
rect 590142 709082 590698 709638
rect 589182 708122 589738 708678
rect 588222 707162 588778 707718
rect 581546 706202 582102 706758
rect 570986 680058 571542 680614
rect 570986 644058 571542 644614
rect 570986 608058 571542 608614
rect 570986 572058 571542 572614
rect 570986 536058 571542 536614
rect 570986 500058 571542 500614
rect 570986 464058 571542 464614
rect 570986 428058 571542 428614
rect 570986 392058 571542 392614
rect 570986 356058 571542 356614
rect 570986 320058 571542 320614
rect 570986 284058 571542 284614
rect 570986 248058 571542 248614
rect 570986 212058 571542 212614
rect 570986 176058 571542 176614
rect 570986 140058 571542 140614
rect 570986 104058 571542 104614
rect 570986 68058 571542 68614
rect 570986 32058 571542 32614
rect 552986 -6662 553542 -6106
rect 577826 704282 578382 704838
rect 577826 686898 578382 687454
rect 577826 650898 578382 651454
rect 577826 614898 578382 615454
rect 577826 578898 578382 579454
rect 577826 542898 578382 543454
rect 577826 506898 578382 507454
rect 577826 470898 578382 471454
rect 577826 434898 578382 435454
rect 577826 398898 578382 399454
rect 577826 362898 578382 363454
rect 577826 326898 578382 327454
rect 577826 290898 578382 291454
rect 577826 254898 578382 255454
rect 577826 218898 578382 219454
rect 577826 182898 578382 183454
rect 577826 146898 578382 147454
rect 577826 110898 578382 111454
rect 577826 74898 578382 75454
rect 577826 38898 578382 39454
rect 577826 2898 578382 3454
rect 577826 -902 578382 -346
rect 587262 706202 587818 706758
rect 586302 705242 586858 705798
rect 581546 690618 582102 691174
rect 581546 654618 582102 655174
rect 581546 618618 582102 619174
rect 581546 582618 582102 583174
rect 581546 546618 582102 547174
rect 581546 510618 582102 511174
rect 581546 474618 582102 475174
rect 581546 438618 582102 439174
rect 581546 402618 582102 403174
rect 581546 366618 582102 367174
rect 581546 330618 582102 331174
rect 581546 294618 582102 295174
rect 581546 258618 582102 259174
rect 581546 222618 582102 223174
rect 581546 186618 582102 187174
rect 581546 150618 582102 151174
rect 581546 114618 582102 115174
rect 581546 78618 582102 79174
rect 581546 42618 582102 43174
rect 581546 6618 582102 7174
rect 585342 704282 585898 704838
rect 585342 686898 585898 687454
rect 585342 650898 585898 651454
rect 585342 614898 585898 615454
rect 585342 578898 585898 579454
rect 585342 542898 585898 543454
rect 585342 506898 585898 507454
rect 585342 470898 585898 471454
rect 585342 434898 585898 435454
rect 585342 398898 585898 399454
rect 585342 362898 585898 363454
rect 585342 326898 585898 327454
rect 585342 290898 585898 291454
rect 585342 254898 585898 255454
rect 585342 218898 585898 219454
rect 585342 182898 585898 183454
rect 585342 146898 585898 147454
rect 585342 110898 585898 111454
rect 585342 74898 585898 75454
rect 585342 38898 585898 39454
rect 585342 2898 585898 3454
rect 585342 -902 585898 -346
rect 586302 668898 586858 669454
rect 586302 632898 586858 633454
rect 586302 596898 586858 597454
rect 586302 560898 586858 561454
rect 586302 524898 586858 525454
rect 586302 488898 586858 489454
rect 586302 452898 586858 453454
rect 586302 416898 586858 417454
rect 586302 380898 586858 381454
rect 586302 344898 586858 345454
rect 586302 308898 586858 309454
rect 586302 272898 586858 273454
rect 586302 236898 586858 237454
rect 586302 200898 586858 201454
rect 586302 164898 586858 165454
rect 586302 128898 586858 129454
rect 586302 92898 586858 93454
rect 586302 56898 586858 57454
rect 586302 20898 586858 21454
rect 586302 -1862 586858 -1306
rect 587262 690618 587818 691174
rect 587262 654618 587818 655174
rect 587262 618618 587818 619174
rect 587262 582618 587818 583174
rect 587262 546618 587818 547174
rect 587262 510618 587818 511174
rect 587262 474618 587818 475174
rect 587262 438618 587818 439174
rect 587262 402618 587818 403174
rect 587262 366618 587818 367174
rect 587262 330618 587818 331174
rect 587262 294618 587818 295174
rect 587262 258618 587818 259174
rect 587262 222618 587818 223174
rect 587262 186618 587818 187174
rect 587262 150618 587818 151174
rect 587262 114618 587818 115174
rect 587262 78618 587818 79174
rect 587262 42618 587818 43174
rect 587262 6618 587818 7174
rect 581546 -2822 582102 -2266
rect 587262 -2822 587818 -2266
rect 588222 672618 588778 673174
rect 588222 636618 588778 637174
rect 588222 600618 588778 601174
rect 588222 564618 588778 565174
rect 588222 528618 588778 529174
rect 588222 492618 588778 493174
rect 588222 456618 588778 457174
rect 588222 420618 588778 421174
rect 588222 384618 588778 385174
rect 588222 348618 588778 349174
rect 588222 312618 588778 313174
rect 588222 276618 588778 277174
rect 588222 240618 588778 241174
rect 588222 204618 588778 205174
rect 588222 168618 588778 169174
rect 588222 132618 588778 133174
rect 588222 96618 588778 97174
rect 588222 60618 588778 61174
rect 588222 24618 588778 25174
rect 588222 -3782 588778 -3226
rect 589182 694338 589738 694894
rect 589182 658338 589738 658894
rect 589182 622338 589738 622894
rect 589182 586338 589738 586894
rect 589182 550338 589738 550894
rect 589182 514338 589738 514894
rect 589182 478338 589738 478894
rect 589182 442338 589738 442894
rect 589182 406338 589738 406894
rect 589182 370338 589738 370894
rect 589182 334338 589738 334894
rect 589182 298338 589738 298894
rect 589182 262338 589738 262894
rect 589182 226338 589738 226894
rect 589182 190338 589738 190894
rect 589182 154338 589738 154894
rect 589182 118338 589738 118894
rect 589182 82338 589738 82894
rect 589182 46338 589738 46894
rect 589182 10338 589738 10894
rect 589182 -4742 589738 -4186
rect 590142 676338 590698 676894
rect 590142 640338 590698 640894
rect 590142 604338 590698 604894
rect 590142 568338 590698 568894
rect 590142 532338 590698 532894
rect 590142 496338 590698 496894
rect 590142 460338 590698 460894
rect 590142 424338 590698 424894
rect 590142 388338 590698 388894
rect 590142 352338 590698 352894
rect 590142 316338 590698 316894
rect 590142 280338 590698 280894
rect 590142 244338 590698 244894
rect 590142 208338 590698 208894
rect 590142 172338 590698 172894
rect 590142 136338 590698 136894
rect 590142 100338 590698 100894
rect 590142 64338 590698 64894
rect 590142 28338 590698 28894
rect 590142 -5702 590698 -5146
rect 591102 698058 591658 698614
rect 591102 662058 591658 662614
rect 591102 626058 591658 626614
rect 591102 590058 591658 590614
rect 591102 554058 591658 554614
rect 591102 518058 591658 518614
rect 591102 482058 591658 482614
rect 591102 446058 591658 446614
rect 591102 410058 591658 410614
rect 591102 374058 591658 374614
rect 591102 338058 591658 338614
rect 591102 302058 591658 302614
rect 591102 266058 591658 266614
rect 591102 230058 591658 230614
rect 591102 194058 591658 194614
rect 591102 158058 591658 158614
rect 591102 122058 591658 122614
rect 591102 86058 591658 86614
rect 591102 50058 591658 50614
rect 591102 14058 591658 14614
rect 591102 -6662 591658 -6106
rect 592062 680058 592618 680614
rect 592062 644058 592618 644614
rect 592062 608058 592618 608614
rect 592062 572058 592618 572614
rect 592062 536058 592618 536614
rect 592062 500058 592618 500614
rect 592062 464058 592618 464614
rect 592062 428058 592618 428614
rect 592062 392058 592618 392614
rect 592062 356058 592618 356614
rect 592062 320058 592618 320614
rect 592062 284058 592618 284614
rect 592062 248058 592618 248614
rect 592062 212058 592618 212614
rect 592062 176058 592618 176614
rect 592062 140058 592618 140614
rect 592062 104058 592618 104614
rect 592062 68058 592618 68614
rect 592062 32058 592618 32614
rect 570986 -7622 571542 -7066
rect 592062 -7622 592618 -7066
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711002 -8694 711558
rect -8138 711002 30986 711558
rect 31542 711002 66986 711558
rect 67542 711002 102986 711558
rect 103542 711002 138986 711558
rect 139542 711002 174986 711558
rect 175542 711002 210986 711558
rect 211542 711002 246986 711558
rect 247542 711002 282986 711558
rect 283542 711002 318986 711558
rect 319542 711002 354986 711558
rect 355542 711002 390986 711558
rect 391542 711002 426986 711558
rect 427542 711002 462986 711558
rect 463542 711002 498986 711558
rect 499542 711002 534986 711558
rect 535542 711002 570986 711558
rect 571542 711002 592062 711558
rect 592618 711002 592650 711558
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710042 -7734 710598
rect -7178 710042 12986 710598
rect 13542 710042 48986 710598
rect 49542 710042 84986 710598
rect 85542 710042 120986 710598
rect 121542 710042 156986 710598
rect 157542 710042 192986 710598
rect 193542 710042 228986 710598
rect 229542 710042 264986 710598
rect 265542 710042 300986 710598
rect 301542 710042 336986 710598
rect 337542 710042 372986 710598
rect 373542 710042 408986 710598
rect 409542 710042 444986 710598
rect 445542 710042 480986 710598
rect 481542 710042 516986 710598
rect 517542 710042 552986 710598
rect 553542 710042 591102 710598
rect 591658 710042 591690 710598
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709082 -6774 709638
rect -6218 709082 27266 709638
rect 27822 709082 63266 709638
rect 63822 709082 99266 709638
rect 99822 709082 135266 709638
rect 135822 709082 171266 709638
rect 171822 709082 207266 709638
rect 207822 709082 243266 709638
rect 243822 709082 279266 709638
rect 279822 709082 315266 709638
rect 315822 709082 351266 709638
rect 351822 709082 387266 709638
rect 387822 709082 423266 709638
rect 423822 709082 459266 709638
rect 459822 709082 495266 709638
rect 495822 709082 531266 709638
rect 531822 709082 567266 709638
rect 567822 709082 590142 709638
rect 590698 709082 590730 709638
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708122 -5814 708678
rect -5258 708122 9266 708678
rect 9822 708122 45266 708678
rect 45822 708122 81266 708678
rect 81822 708122 117266 708678
rect 117822 708122 153266 708678
rect 153822 708122 189266 708678
rect 189822 708122 225266 708678
rect 225822 708122 261266 708678
rect 261822 708122 297266 708678
rect 297822 708122 333266 708678
rect 333822 708122 369266 708678
rect 369822 708122 405266 708678
rect 405822 708122 441266 708678
rect 441822 708122 477266 708678
rect 477822 708122 513266 708678
rect 513822 708122 549266 708678
rect 549822 708122 589182 708678
rect 589738 708122 589770 708678
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707162 -4854 707718
rect -4298 707162 23546 707718
rect 24102 707162 59546 707718
rect 60102 707162 95546 707718
rect 96102 707162 131546 707718
rect 132102 707162 167546 707718
rect 168102 707162 203546 707718
rect 204102 707162 239546 707718
rect 240102 707162 275546 707718
rect 276102 707162 311546 707718
rect 312102 707162 347546 707718
rect 348102 707162 383546 707718
rect 384102 707162 419546 707718
rect 420102 707162 455546 707718
rect 456102 707162 491546 707718
rect 492102 707162 527546 707718
rect 528102 707162 563546 707718
rect 564102 707162 588222 707718
rect 588778 707162 588810 707718
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706202 -3894 706758
rect -3338 706202 5546 706758
rect 6102 706202 41546 706758
rect 42102 706202 77546 706758
rect 78102 706202 113546 706758
rect 114102 706202 149546 706758
rect 150102 706202 185546 706758
rect 186102 706202 221546 706758
rect 222102 706202 257546 706758
rect 258102 706202 293546 706758
rect 294102 706202 329546 706758
rect 330102 706202 365546 706758
rect 366102 706202 401546 706758
rect 402102 706202 437546 706758
rect 438102 706202 473546 706758
rect 474102 706202 509546 706758
rect 510102 706202 545546 706758
rect 546102 706202 581546 706758
rect 582102 706202 587262 706758
rect 587818 706202 587850 706758
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705242 -2934 705798
rect -2378 705242 19826 705798
rect 20382 705242 55826 705798
rect 56382 705242 91826 705798
rect 92382 705242 127826 705798
rect 128382 705242 163826 705798
rect 164382 705242 199826 705798
rect 200382 705242 235826 705798
rect 236382 705242 271826 705798
rect 272382 705242 307826 705798
rect 308382 705242 343826 705798
rect 344382 705242 379826 705798
rect 380382 705242 415826 705798
rect 416382 705242 451826 705798
rect 452382 705242 487826 705798
rect 488382 705242 523826 705798
rect 524382 705242 559826 705798
rect 560382 705242 586302 705798
rect 586858 705242 586890 705798
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704282 -1974 704838
rect -1418 704282 1826 704838
rect 2382 704282 37826 704838
rect 38382 704282 73826 704838
rect 74382 704282 109826 704838
rect 110382 704282 145826 704838
rect 146382 704282 181826 704838
rect 182382 704282 217826 704838
rect 218382 704282 253826 704838
rect 254382 704282 289826 704838
rect 290382 704282 325826 704838
rect 326382 704282 361826 704838
rect 362382 704282 397826 704838
rect 398382 704282 433826 704838
rect 434382 704282 469826 704838
rect 470382 704282 505826 704838
rect 506382 704282 541826 704838
rect 542382 704282 577826 704838
rect 578382 704282 585342 704838
rect 585898 704282 585930 704838
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698058 -7734 698614
rect -7178 698058 12986 698614
rect 13542 698058 48986 698614
rect 49542 698058 84986 698614
rect 85542 698058 120986 698614
rect 121542 698058 156986 698614
rect 157542 698058 192986 698614
rect 193542 698058 228986 698614
rect 229542 698058 264986 698614
rect 265542 698058 300986 698614
rect 301542 698058 336986 698614
rect 337542 698058 372986 698614
rect 373542 698058 408986 698614
rect 409542 698058 444986 698614
rect 445542 698058 480986 698614
rect 481542 698058 516986 698614
rect 517542 698058 552986 698614
rect 553542 698058 591102 698614
rect 591658 698058 592650 698614
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694338 -5814 694894
rect -5258 694338 9266 694894
rect 9822 694338 45266 694894
rect 45822 694338 81266 694894
rect 81822 694338 117266 694894
rect 117822 694338 153266 694894
rect 153822 694338 189266 694894
rect 189822 694338 225266 694894
rect 225822 694338 261266 694894
rect 261822 694338 297266 694894
rect 297822 694338 333266 694894
rect 333822 694338 369266 694894
rect 369822 694338 405266 694894
rect 405822 694338 441266 694894
rect 441822 694338 477266 694894
rect 477822 694338 513266 694894
rect 513822 694338 549266 694894
rect 549822 694338 589182 694894
rect 589738 694338 590730 694894
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690618 -3894 691174
rect -3338 690618 5546 691174
rect 6102 690618 41546 691174
rect 42102 690618 77546 691174
rect 78102 690618 113546 691174
rect 114102 690618 149546 691174
rect 150102 690618 185546 691174
rect 186102 690618 221546 691174
rect 222102 690618 257546 691174
rect 258102 690618 293546 691174
rect 294102 690618 329546 691174
rect 330102 690618 365546 691174
rect 366102 690618 401546 691174
rect 402102 690618 437546 691174
rect 438102 690618 473546 691174
rect 474102 690618 509546 691174
rect 510102 690618 545546 691174
rect 546102 690618 581546 691174
rect 582102 690618 587262 691174
rect 587818 690618 588810 691174
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 686898 -1974 687454
rect -1418 686898 1826 687454
rect 2382 686898 37826 687454
rect 38382 686898 73826 687454
rect 74382 686898 109826 687454
rect 110382 686898 145826 687454
rect 146382 686898 181826 687454
rect 182382 686898 217826 687454
rect 218382 686898 253826 687454
rect 254382 686898 289826 687454
rect 290382 686898 325826 687454
rect 326382 686898 361826 687454
rect 362382 686898 397826 687454
rect 398382 686898 433826 687454
rect 434382 686898 469826 687454
rect 470382 686898 505826 687454
rect 506382 686898 541826 687454
rect 542382 686898 577826 687454
rect 578382 686898 585342 687454
rect 585898 686898 586890 687454
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680058 -8694 680614
rect -8138 680058 30986 680614
rect 31542 680058 66986 680614
rect 67542 680058 102986 680614
rect 103542 680058 138986 680614
rect 139542 680058 174986 680614
rect 175542 680058 210986 680614
rect 211542 680058 246986 680614
rect 247542 680058 282986 680614
rect 283542 680058 318986 680614
rect 319542 680058 354986 680614
rect 355542 680058 390986 680614
rect 391542 680058 426986 680614
rect 427542 680058 462986 680614
rect 463542 680058 498986 680614
rect 499542 680058 534986 680614
rect 535542 680058 570986 680614
rect 571542 680058 592062 680614
rect 592618 680058 592650 680614
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676338 -6774 676894
rect -6218 676338 27266 676894
rect 27822 676338 63266 676894
rect 63822 676338 99266 676894
rect 99822 676338 135266 676894
rect 135822 676338 171266 676894
rect 171822 676338 207266 676894
rect 207822 676338 243266 676894
rect 243822 676338 279266 676894
rect 279822 676338 315266 676894
rect 315822 676338 351266 676894
rect 351822 676338 387266 676894
rect 387822 676338 423266 676894
rect 423822 676338 459266 676894
rect 459822 676338 495266 676894
rect 495822 676338 531266 676894
rect 531822 676338 567266 676894
rect 567822 676338 590142 676894
rect 590698 676338 590730 676894
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672618 -4854 673174
rect -4298 672618 23546 673174
rect 24102 672618 59546 673174
rect 60102 672618 95546 673174
rect 96102 672618 131546 673174
rect 132102 672618 167546 673174
rect 168102 672618 203546 673174
rect 204102 672618 239546 673174
rect 240102 672618 275546 673174
rect 276102 672618 311546 673174
rect 312102 672618 347546 673174
rect 348102 672618 383546 673174
rect 384102 672618 419546 673174
rect 420102 672618 455546 673174
rect 456102 672618 491546 673174
rect 492102 672618 527546 673174
rect 528102 672618 563546 673174
rect 564102 672618 588222 673174
rect 588778 672618 588810 673174
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 668898 -2934 669454
rect -2378 668898 19826 669454
rect 20382 668898 55826 669454
rect 56382 668898 91826 669454
rect 92382 668898 127826 669454
rect 128382 668898 163826 669454
rect 164382 668898 199826 669454
rect 200382 668898 235826 669454
rect 236382 668898 271826 669454
rect 272382 668898 307826 669454
rect 308382 668898 343826 669454
rect 344382 668898 379826 669454
rect 380382 668898 415826 669454
rect 416382 668898 451826 669454
rect 452382 668898 487826 669454
rect 488382 668898 523826 669454
rect 524382 668898 559826 669454
rect 560382 668898 586302 669454
rect 586858 668898 586890 669454
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662058 -7734 662614
rect -7178 662058 12986 662614
rect 13542 662058 48986 662614
rect 49542 662058 84986 662614
rect 85542 662058 120986 662614
rect 121542 662058 156986 662614
rect 157542 662058 192986 662614
rect 193542 662058 228986 662614
rect 229542 662058 264986 662614
rect 265542 662058 300986 662614
rect 301542 662058 336986 662614
rect 337542 662058 372986 662614
rect 373542 662058 408986 662614
rect 409542 662058 444986 662614
rect 445542 662058 480986 662614
rect 481542 662058 516986 662614
rect 517542 662058 552986 662614
rect 553542 662058 591102 662614
rect 591658 662058 592650 662614
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658338 -5814 658894
rect -5258 658338 9266 658894
rect 9822 658338 45266 658894
rect 45822 658338 81266 658894
rect 81822 658338 117266 658894
rect 117822 658338 153266 658894
rect 153822 658338 189266 658894
rect 189822 658338 225266 658894
rect 225822 658338 261266 658894
rect 261822 658338 297266 658894
rect 297822 658338 333266 658894
rect 333822 658338 369266 658894
rect 369822 658338 405266 658894
rect 405822 658338 441266 658894
rect 441822 658338 477266 658894
rect 477822 658338 513266 658894
rect 513822 658338 549266 658894
rect 549822 658338 589182 658894
rect 589738 658338 590730 658894
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654618 -3894 655174
rect -3338 654618 5546 655174
rect 6102 654618 41546 655174
rect 42102 654618 77546 655174
rect 78102 654618 113546 655174
rect 114102 654618 149546 655174
rect 150102 654618 185546 655174
rect 186102 654618 221546 655174
rect 222102 654618 257546 655174
rect 258102 654618 293546 655174
rect 294102 654618 329546 655174
rect 330102 654618 365546 655174
rect 366102 654618 401546 655174
rect 402102 654618 437546 655174
rect 438102 654618 473546 655174
rect 474102 654618 509546 655174
rect 510102 654618 545546 655174
rect 546102 654618 581546 655174
rect 582102 654618 587262 655174
rect 587818 654618 588810 655174
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 650898 -1974 651454
rect -1418 650898 1826 651454
rect 2382 650898 37826 651454
rect 38382 650898 73826 651454
rect 74382 650898 109826 651454
rect 110382 650898 145826 651454
rect 146382 650898 181826 651454
rect 182382 650898 217826 651454
rect 218382 650898 253826 651454
rect 254382 650898 289826 651454
rect 290382 650898 325826 651454
rect 326382 650898 361826 651454
rect 362382 650898 397826 651454
rect 398382 650898 433826 651454
rect 434382 650898 469826 651454
rect 470382 650898 505826 651454
rect 506382 650898 541826 651454
rect 542382 650898 577826 651454
rect 578382 650898 585342 651454
rect 585898 650898 586890 651454
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644058 -8694 644614
rect -8138 644058 30986 644614
rect 31542 644058 66986 644614
rect 67542 644058 102986 644614
rect 103542 644058 138986 644614
rect 139542 644058 174986 644614
rect 175542 644058 210986 644614
rect 211542 644058 246986 644614
rect 247542 644058 282986 644614
rect 283542 644058 318986 644614
rect 319542 644058 354986 644614
rect 355542 644058 390986 644614
rect 391542 644058 426986 644614
rect 427542 644058 462986 644614
rect 463542 644058 498986 644614
rect 499542 644058 534986 644614
rect 535542 644058 570986 644614
rect 571542 644058 592062 644614
rect 592618 644058 592650 644614
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640338 -6774 640894
rect -6218 640338 27266 640894
rect 27822 640338 63266 640894
rect 63822 640338 99266 640894
rect 99822 640338 135266 640894
rect 135822 640338 171266 640894
rect 171822 640338 207266 640894
rect 207822 640338 243266 640894
rect 243822 640338 279266 640894
rect 279822 640338 315266 640894
rect 315822 640338 351266 640894
rect 351822 640338 387266 640894
rect 387822 640338 423266 640894
rect 423822 640338 459266 640894
rect 459822 640338 495266 640894
rect 495822 640338 531266 640894
rect 531822 640338 567266 640894
rect 567822 640338 590142 640894
rect 590698 640338 590730 640894
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636618 -4854 637174
rect -4298 636618 23546 637174
rect 24102 636618 59546 637174
rect 60102 636618 95546 637174
rect 96102 636618 131546 637174
rect 132102 636618 167546 637174
rect 168102 636618 203546 637174
rect 204102 636618 239546 637174
rect 240102 636618 275546 637174
rect 276102 636618 311546 637174
rect 312102 636618 347546 637174
rect 348102 636618 383546 637174
rect 384102 636618 419546 637174
rect 420102 636618 455546 637174
rect 456102 636618 491546 637174
rect 492102 636618 527546 637174
rect 528102 636618 563546 637174
rect 564102 636618 588222 637174
rect 588778 636618 588810 637174
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 632898 -2934 633454
rect -2378 632898 19826 633454
rect 20382 632898 55826 633454
rect 56382 632898 91826 633454
rect 92382 632898 127826 633454
rect 128382 632898 163826 633454
rect 164382 632898 199826 633454
rect 200382 632898 235826 633454
rect 236382 632898 271826 633454
rect 272382 632898 307826 633454
rect 308382 632898 343826 633454
rect 344382 632898 379826 633454
rect 380382 632898 415826 633454
rect 416382 632898 451826 633454
rect 452382 632898 487826 633454
rect 488382 632898 523826 633454
rect 524382 632898 559826 633454
rect 560382 632898 586302 633454
rect 586858 632898 586890 633454
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626058 -7734 626614
rect -7178 626058 12986 626614
rect 13542 626058 48986 626614
rect 49542 626058 84986 626614
rect 85542 626058 120986 626614
rect 121542 626058 156986 626614
rect 157542 626058 192986 626614
rect 193542 626058 228986 626614
rect 229542 626058 264986 626614
rect 265542 626058 300986 626614
rect 301542 626058 336986 626614
rect 337542 626058 372986 626614
rect 373542 626058 408986 626614
rect 409542 626058 444986 626614
rect 445542 626058 480986 626614
rect 481542 626058 516986 626614
rect 517542 626058 552986 626614
rect 553542 626058 591102 626614
rect 591658 626058 592650 626614
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622338 -5814 622894
rect -5258 622338 9266 622894
rect 9822 622338 45266 622894
rect 45822 622338 81266 622894
rect 81822 622338 117266 622894
rect 117822 622338 153266 622894
rect 153822 622338 189266 622894
rect 189822 622338 225266 622894
rect 225822 622338 261266 622894
rect 261822 622338 297266 622894
rect 297822 622338 333266 622894
rect 333822 622338 369266 622894
rect 369822 622338 405266 622894
rect 405822 622338 441266 622894
rect 441822 622338 477266 622894
rect 477822 622338 513266 622894
rect 513822 622338 549266 622894
rect 549822 622338 589182 622894
rect 589738 622338 590730 622894
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618618 -3894 619174
rect -3338 618618 5546 619174
rect 6102 618618 41546 619174
rect 42102 618618 77546 619174
rect 78102 618618 113546 619174
rect 114102 618618 149546 619174
rect 150102 618618 185546 619174
rect 186102 618618 221546 619174
rect 222102 618618 257546 619174
rect 258102 618618 293546 619174
rect 294102 618618 329546 619174
rect 330102 618618 365546 619174
rect 366102 618618 401546 619174
rect 402102 618618 437546 619174
rect 438102 618618 473546 619174
rect 474102 618618 509546 619174
rect 510102 618618 545546 619174
rect 546102 618618 581546 619174
rect 582102 618618 587262 619174
rect 587818 618618 588810 619174
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 614898 -1974 615454
rect -1418 614898 1826 615454
rect 2382 614898 37826 615454
rect 38382 614898 73826 615454
rect 74382 614898 109826 615454
rect 110382 614898 145826 615454
rect 146382 614898 181826 615454
rect 182382 614898 217826 615454
rect 218382 614898 253826 615454
rect 254382 614898 289826 615454
rect 290382 614898 325826 615454
rect 326382 614898 361826 615454
rect 362382 614898 397826 615454
rect 398382 614898 433826 615454
rect 434382 614898 469826 615454
rect 470382 614898 505826 615454
rect 506382 614898 541826 615454
rect 542382 614898 577826 615454
rect 578382 614898 585342 615454
rect 585898 614898 586890 615454
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608058 -8694 608614
rect -8138 608058 30986 608614
rect 31542 608058 66986 608614
rect 67542 608058 102986 608614
rect 103542 608058 138986 608614
rect 139542 608058 174986 608614
rect 175542 608058 210986 608614
rect 211542 608058 246986 608614
rect 247542 608058 282986 608614
rect 283542 608058 318986 608614
rect 319542 608058 354986 608614
rect 355542 608058 390986 608614
rect 391542 608058 426986 608614
rect 427542 608058 462986 608614
rect 463542 608058 498986 608614
rect 499542 608058 534986 608614
rect 535542 608058 570986 608614
rect 571542 608058 592062 608614
rect 592618 608058 592650 608614
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604338 -6774 604894
rect -6218 604338 27266 604894
rect 27822 604338 63266 604894
rect 63822 604338 99266 604894
rect 99822 604338 135266 604894
rect 135822 604338 171266 604894
rect 171822 604338 207266 604894
rect 207822 604338 243266 604894
rect 243822 604338 279266 604894
rect 279822 604338 315266 604894
rect 315822 604338 351266 604894
rect 351822 604338 387266 604894
rect 387822 604338 423266 604894
rect 423822 604338 459266 604894
rect 459822 604338 495266 604894
rect 495822 604338 531266 604894
rect 531822 604338 567266 604894
rect 567822 604338 590142 604894
rect 590698 604338 590730 604894
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600618 -4854 601174
rect -4298 600618 23546 601174
rect 24102 600618 59546 601174
rect 60102 600618 95546 601174
rect 96102 600618 131546 601174
rect 132102 600618 167546 601174
rect 168102 600618 203546 601174
rect 204102 600618 239546 601174
rect 240102 600618 275546 601174
rect 276102 600618 311546 601174
rect 312102 600618 347546 601174
rect 348102 600618 383546 601174
rect 384102 600618 419546 601174
rect 420102 600618 455546 601174
rect 456102 600618 491546 601174
rect 492102 600618 527546 601174
rect 528102 600618 563546 601174
rect 564102 600618 588222 601174
rect 588778 600618 588810 601174
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 596898 -2934 597454
rect -2378 596898 19826 597454
rect 20382 596898 55826 597454
rect 56382 596898 91826 597454
rect 92382 596898 127826 597454
rect 128382 596898 163826 597454
rect 164382 596898 199826 597454
rect 200382 596898 235826 597454
rect 236382 596898 271826 597454
rect 272382 596898 307826 597454
rect 308382 596898 343826 597454
rect 344382 596898 379826 597454
rect 380382 596898 415826 597454
rect 416382 596898 451826 597454
rect 452382 596898 487826 597454
rect 488382 596898 523826 597454
rect 524382 596898 559826 597454
rect 560382 596898 586302 597454
rect 586858 596898 586890 597454
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590058 -7734 590614
rect -7178 590058 12986 590614
rect 13542 590058 48986 590614
rect 49542 590058 84986 590614
rect 85542 590058 120986 590614
rect 121542 590058 156986 590614
rect 157542 590058 192986 590614
rect 193542 590058 228986 590614
rect 229542 590058 264986 590614
rect 265542 590058 300986 590614
rect 301542 590058 336986 590614
rect 337542 590058 372986 590614
rect 373542 590058 408986 590614
rect 409542 590058 444986 590614
rect 445542 590058 480986 590614
rect 481542 590058 516986 590614
rect 517542 590058 552986 590614
rect 553542 590058 591102 590614
rect 591658 590058 592650 590614
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586338 -5814 586894
rect -5258 586338 9266 586894
rect 9822 586338 45266 586894
rect 45822 586338 81266 586894
rect 81822 586338 117266 586894
rect 117822 586338 153266 586894
rect 153822 586338 189266 586894
rect 189822 586338 225266 586894
rect 225822 586338 261266 586894
rect 261822 586338 297266 586894
rect 297822 586338 333266 586894
rect 333822 586338 369266 586894
rect 369822 586338 405266 586894
rect 405822 586338 441266 586894
rect 441822 586338 477266 586894
rect 477822 586338 513266 586894
rect 513822 586338 549266 586894
rect 549822 586338 589182 586894
rect 589738 586338 590730 586894
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582618 -3894 583174
rect -3338 582618 5546 583174
rect 6102 582618 41546 583174
rect 42102 582618 77546 583174
rect 78102 582618 113546 583174
rect 114102 582618 149546 583174
rect 150102 582618 185546 583174
rect 186102 582618 221546 583174
rect 222102 582618 257546 583174
rect 258102 582618 293546 583174
rect 294102 582618 329546 583174
rect 330102 582618 365546 583174
rect 366102 582618 401546 583174
rect 402102 582618 437546 583174
rect 438102 582618 473546 583174
rect 474102 582618 509546 583174
rect 510102 582618 545546 583174
rect 546102 582618 581546 583174
rect 582102 582618 587262 583174
rect 587818 582618 588810 583174
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 578898 -1974 579454
rect -1418 578898 1826 579454
rect 2382 578898 37826 579454
rect 38382 578898 73826 579454
rect 74382 578898 109826 579454
rect 110382 578898 145826 579454
rect 146382 578898 181826 579454
rect 182382 578898 217826 579454
rect 218382 578898 253826 579454
rect 254382 578898 289826 579454
rect 290382 578898 325826 579454
rect 326382 578898 361826 579454
rect 362382 578898 397826 579454
rect 398382 578898 433826 579454
rect 434382 578898 469826 579454
rect 470382 578898 505826 579454
rect 506382 578898 541826 579454
rect 542382 578898 577826 579454
rect 578382 578898 585342 579454
rect 585898 578898 586890 579454
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572058 -8694 572614
rect -8138 572058 30986 572614
rect 31542 572058 66986 572614
rect 67542 572058 102986 572614
rect 103542 572058 138986 572614
rect 139542 572058 174986 572614
rect 175542 572058 210986 572614
rect 211542 572058 246986 572614
rect 247542 572058 282986 572614
rect 283542 572058 318986 572614
rect 319542 572058 354986 572614
rect 355542 572058 390986 572614
rect 391542 572058 426986 572614
rect 427542 572058 462986 572614
rect 463542 572058 498986 572614
rect 499542 572058 534986 572614
rect 535542 572058 570986 572614
rect 571542 572058 592062 572614
rect 592618 572058 592650 572614
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568338 -6774 568894
rect -6218 568338 27266 568894
rect 27822 568338 63266 568894
rect 63822 568338 99266 568894
rect 99822 568338 135266 568894
rect 135822 568338 171266 568894
rect 171822 568338 207266 568894
rect 207822 568338 243266 568894
rect 243822 568338 279266 568894
rect 279822 568338 315266 568894
rect 315822 568338 351266 568894
rect 351822 568338 387266 568894
rect 387822 568338 423266 568894
rect 423822 568338 459266 568894
rect 459822 568338 495266 568894
rect 495822 568338 531266 568894
rect 531822 568338 567266 568894
rect 567822 568338 590142 568894
rect 590698 568338 590730 568894
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564618 -4854 565174
rect -4298 564618 23546 565174
rect 24102 564618 59546 565174
rect 60102 564618 95546 565174
rect 96102 564618 131546 565174
rect 132102 564618 167546 565174
rect 168102 564618 203546 565174
rect 204102 564618 239546 565174
rect 240102 564618 275546 565174
rect 276102 564618 311546 565174
rect 312102 564618 347546 565174
rect 348102 564618 383546 565174
rect 384102 564618 419546 565174
rect 420102 564618 455546 565174
rect 456102 564618 491546 565174
rect 492102 564618 527546 565174
rect 528102 564618 563546 565174
rect 564102 564618 588222 565174
rect 588778 564618 588810 565174
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 560898 -2934 561454
rect -2378 560898 19826 561454
rect 20382 560898 55826 561454
rect 56382 560898 91826 561454
rect 92382 560898 127826 561454
rect 128382 560898 163826 561454
rect 164382 560898 199826 561454
rect 200382 560898 235826 561454
rect 236382 560898 271826 561454
rect 272382 560898 307826 561454
rect 308382 560898 343826 561454
rect 344382 560898 379826 561454
rect 380382 560898 415826 561454
rect 416382 560898 451826 561454
rect 452382 560898 487826 561454
rect 488382 560898 523826 561454
rect 524382 560898 559826 561454
rect 560382 560898 586302 561454
rect 586858 560898 586890 561454
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554058 -7734 554614
rect -7178 554058 12986 554614
rect 13542 554058 48986 554614
rect 49542 554058 84986 554614
rect 85542 554058 120986 554614
rect 121542 554058 156986 554614
rect 157542 554058 192986 554614
rect 193542 554058 228986 554614
rect 229542 554058 264986 554614
rect 265542 554058 300986 554614
rect 301542 554058 336986 554614
rect 337542 554058 372986 554614
rect 373542 554058 408986 554614
rect 409542 554058 444986 554614
rect 445542 554058 480986 554614
rect 481542 554058 516986 554614
rect 517542 554058 552986 554614
rect 553542 554058 591102 554614
rect 591658 554058 592650 554614
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550338 -5814 550894
rect -5258 550338 9266 550894
rect 9822 550338 45266 550894
rect 45822 550338 81266 550894
rect 81822 550338 117266 550894
rect 117822 550338 153266 550894
rect 153822 550338 189266 550894
rect 189822 550338 225266 550894
rect 225822 550338 261266 550894
rect 261822 550338 297266 550894
rect 297822 550338 333266 550894
rect 333822 550338 369266 550894
rect 369822 550338 405266 550894
rect 405822 550338 441266 550894
rect 441822 550338 477266 550894
rect 477822 550338 513266 550894
rect 513822 550338 549266 550894
rect 549822 550338 589182 550894
rect 589738 550338 590730 550894
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546618 -3894 547174
rect -3338 546618 5546 547174
rect 6102 546618 41546 547174
rect 42102 546618 77546 547174
rect 78102 546618 113546 547174
rect 114102 546618 149546 547174
rect 150102 546618 185546 547174
rect 186102 546618 221546 547174
rect 222102 546618 257546 547174
rect 258102 546618 293546 547174
rect 294102 546618 329546 547174
rect 330102 546618 365546 547174
rect 366102 546618 401546 547174
rect 402102 546618 437546 547174
rect 438102 546618 473546 547174
rect 474102 546618 509546 547174
rect 510102 546618 545546 547174
rect 546102 546618 581546 547174
rect 582102 546618 587262 547174
rect 587818 546618 588810 547174
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 542898 -1974 543454
rect -1418 542898 1826 543454
rect 2382 542898 37826 543454
rect 38382 542898 73826 543454
rect 74382 542898 109826 543454
rect 110382 542898 145826 543454
rect 146382 542898 181826 543454
rect 182382 542898 217826 543454
rect 218382 542898 253826 543454
rect 254382 542898 289826 543454
rect 290382 542898 325826 543454
rect 326382 542898 361826 543454
rect 362382 542898 397826 543454
rect 398382 542898 433826 543454
rect 434382 542898 469826 543454
rect 470382 542898 505826 543454
rect 506382 542898 541826 543454
rect 542382 542898 577826 543454
rect 578382 542898 585342 543454
rect 585898 542898 586890 543454
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536058 -8694 536614
rect -8138 536058 30986 536614
rect 31542 536058 66986 536614
rect 67542 536058 102986 536614
rect 103542 536058 138986 536614
rect 139542 536058 174986 536614
rect 175542 536058 210986 536614
rect 211542 536058 246986 536614
rect 247542 536058 282986 536614
rect 283542 536058 318986 536614
rect 319542 536058 354986 536614
rect 355542 536058 390986 536614
rect 391542 536058 426986 536614
rect 427542 536058 462986 536614
rect 463542 536058 498986 536614
rect 499542 536058 534986 536614
rect 535542 536058 570986 536614
rect 571542 536058 592062 536614
rect 592618 536058 592650 536614
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532338 -6774 532894
rect -6218 532338 27266 532894
rect 27822 532338 63266 532894
rect 63822 532338 99266 532894
rect 99822 532338 135266 532894
rect 135822 532338 171266 532894
rect 171822 532338 207266 532894
rect 207822 532338 243266 532894
rect 243822 532338 279266 532894
rect 279822 532338 315266 532894
rect 315822 532338 351266 532894
rect 351822 532338 387266 532894
rect 387822 532338 423266 532894
rect 423822 532338 459266 532894
rect 459822 532338 495266 532894
rect 495822 532338 531266 532894
rect 531822 532338 567266 532894
rect 567822 532338 590142 532894
rect 590698 532338 590730 532894
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528618 -4854 529174
rect -4298 528618 23546 529174
rect 24102 528618 59546 529174
rect 60102 528618 95546 529174
rect 96102 528618 131546 529174
rect 132102 528618 167546 529174
rect 168102 528618 203546 529174
rect 204102 528618 239546 529174
rect 240102 528618 275546 529174
rect 276102 528618 311546 529174
rect 312102 528618 347546 529174
rect 348102 528618 383546 529174
rect 384102 528618 419546 529174
rect 420102 528618 455546 529174
rect 456102 528618 491546 529174
rect 492102 528618 527546 529174
rect 528102 528618 563546 529174
rect 564102 528618 588222 529174
rect 588778 528618 588810 529174
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 524898 -2934 525454
rect -2378 524898 19826 525454
rect 20382 524898 55826 525454
rect 56382 524898 91826 525454
rect 92382 524898 127826 525454
rect 128382 524898 163826 525454
rect 164382 524898 199826 525454
rect 200382 524898 235826 525454
rect 236382 524898 271826 525454
rect 272382 524898 307826 525454
rect 308382 524898 343826 525454
rect 344382 524898 379826 525454
rect 380382 524898 415826 525454
rect 416382 524898 451826 525454
rect 452382 524898 487826 525454
rect 488382 524898 523826 525454
rect 524382 524898 559826 525454
rect 560382 524898 586302 525454
rect 586858 524898 586890 525454
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518058 -7734 518614
rect -7178 518058 12986 518614
rect 13542 518058 48986 518614
rect 49542 518058 84986 518614
rect 85542 518058 120986 518614
rect 121542 518058 156986 518614
rect 157542 518058 192986 518614
rect 193542 518058 228986 518614
rect 229542 518058 264986 518614
rect 265542 518058 300986 518614
rect 301542 518058 336986 518614
rect 337542 518058 372986 518614
rect 373542 518058 408986 518614
rect 409542 518058 444986 518614
rect 445542 518058 480986 518614
rect 481542 518058 516986 518614
rect 517542 518058 552986 518614
rect 553542 518058 591102 518614
rect 591658 518058 592650 518614
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514338 -5814 514894
rect -5258 514338 9266 514894
rect 9822 514338 45266 514894
rect 45822 514338 81266 514894
rect 81822 514338 117266 514894
rect 117822 514338 153266 514894
rect 153822 514338 189266 514894
rect 189822 514338 225266 514894
rect 225822 514338 261266 514894
rect 261822 514338 297266 514894
rect 297822 514338 333266 514894
rect 333822 514338 369266 514894
rect 369822 514338 405266 514894
rect 405822 514338 441266 514894
rect 441822 514338 477266 514894
rect 477822 514338 513266 514894
rect 513822 514338 549266 514894
rect 549822 514338 589182 514894
rect 589738 514338 590730 514894
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510618 -3894 511174
rect -3338 510618 5546 511174
rect 6102 510618 41546 511174
rect 42102 510618 77546 511174
rect 78102 510618 113546 511174
rect 114102 510618 149546 511174
rect 150102 510618 185546 511174
rect 186102 510618 221546 511174
rect 222102 510618 257546 511174
rect 258102 510618 293546 511174
rect 294102 510618 329546 511174
rect 330102 510618 365546 511174
rect 366102 510618 401546 511174
rect 402102 510618 437546 511174
rect 438102 510618 473546 511174
rect 474102 510618 509546 511174
rect 510102 510618 545546 511174
rect 546102 510618 581546 511174
rect 582102 510618 587262 511174
rect 587818 510618 588810 511174
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 506898 -1974 507454
rect -1418 506898 1826 507454
rect 2382 506898 37826 507454
rect 38382 506898 73826 507454
rect 74382 506898 109826 507454
rect 110382 506898 145826 507454
rect 146382 506898 181826 507454
rect 182382 506898 217826 507454
rect 218382 506898 253826 507454
rect 254382 506898 289826 507454
rect 290382 506898 325826 507454
rect 326382 506898 361826 507454
rect 362382 506898 397826 507454
rect 398382 506898 433826 507454
rect 434382 506898 469826 507454
rect 470382 506898 505826 507454
rect 506382 506898 541826 507454
rect 542382 506898 577826 507454
rect 578382 506898 585342 507454
rect 585898 506898 586890 507454
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500058 -8694 500614
rect -8138 500058 30986 500614
rect 31542 500058 66986 500614
rect 67542 500058 102986 500614
rect 103542 500058 138986 500614
rect 139542 500058 174986 500614
rect 175542 500058 210986 500614
rect 211542 500058 246986 500614
rect 247542 500058 282986 500614
rect 283542 500058 318986 500614
rect 319542 500058 354986 500614
rect 355542 500058 390986 500614
rect 391542 500058 426986 500614
rect 427542 500058 462986 500614
rect 463542 500058 498986 500614
rect 499542 500058 534986 500614
rect 535542 500058 570986 500614
rect 571542 500058 592062 500614
rect 592618 500058 592650 500614
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496338 -6774 496894
rect -6218 496338 27266 496894
rect 27822 496338 63266 496894
rect 63822 496338 99266 496894
rect 99822 496338 135266 496894
rect 135822 496338 171266 496894
rect 171822 496338 207266 496894
rect 207822 496338 243266 496894
rect 243822 496338 279266 496894
rect 279822 496338 315266 496894
rect 315822 496338 351266 496894
rect 351822 496338 387266 496894
rect 387822 496338 423266 496894
rect 423822 496338 459266 496894
rect 459822 496338 495266 496894
rect 495822 496338 531266 496894
rect 531822 496338 567266 496894
rect 567822 496338 590142 496894
rect 590698 496338 590730 496894
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492618 -4854 493174
rect -4298 492618 23546 493174
rect 24102 492618 59546 493174
rect 60102 492618 95546 493174
rect 96102 492618 131546 493174
rect 132102 492618 167546 493174
rect 168102 492618 203546 493174
rect 204102 492618 239546 493174
rect 240102 492618 275546 493174
rect 276102 492618 311546 493174
rect 312102 492618 347546 493174
rect 348102 492618 383546 493174
rect 384102 492618 419546 493174
rect 420102 492618 455546 493174
rect 456102 492618 491546 493174
rect 492102 492618 527546 493174
rect 528102 492618 563546 493174
rect 564102 492618 588222 493174
rect 588778 492618 588810 493174
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 488898 -2934 489454
rect -2378 488898 19826 489454
rect 20382 488898 55826 489454
rect 56382 488898 91826 489454
rect 92382 488898 127826 489454
rect 128382 488898 163826 489454
rect 164382 488898 199826 489454
rect 200382 488898 235826 489454
rect 236382 488898 271826 489454
rect 272382 488898 307826 489454
rect 308382 488898 343826 489454
rect 344382 488898 379826 489454
rect 380382 488898 415826 489454
rect 416382 488898 451826 489454
rect 452382 488898 487826 489454
rect 488382 488898 523826 489454
rect 524382 488898 559826 489454
rect 560382 488898 586302 489454
rect 586858 488898 586890 489454
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482058 -7734 482614
rect -7178 482058 12986 482614
rect 13542 482058 48986 482614
rect 49542 482058 84986 482614
rect 85542 482058 120986 482614
rect 121542 482058 156986 482614
rect 157542 482058 192986 482614
rect 193542 482058 228986 482614
rect 229542 482058 264986 482614
rect 265542 482058 300986 482614
rect 301542 482058 336986 482614
rect 337542 482058 372986 482614
rect 373542 482058 408986 482614
rect 409542 482058 444986 482614
rect 445542 482058 480986 482614
rect 481542 482058 516986 482614
rect 517542 482058 552986 482614
rect 553542 482058 591102 482614
rect 591658 482058 592650 482614
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478338 -5814 478894
rect -5258 478338 9266 478894
rect 9822 478338 45266 478894
rect 45822 478338 81266 478894
rect 81822 478338 117266 478894
rect 117822 478338 153266 478894
rect 153822 478338 189266 478894
rect 189822 478338 225266 478894
rect 225822 478338 261266 478894
rect 261822 478338 297266 478894
rect 297822 478338 333266 478894
rect 333822 478338 369266 478894
rect 369822 478338 405266 478894
rect 405822 478338 441266 478894
rect 441822 478338 477266 478894
rect 477822 478338 513266 478894
rect 513822 478338 549266 478894
rect 549822 478338 589182 478894
rect 589738 478338 590730 478894
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474618 -3894 475174
rect -3338 474618 5546 475174
rect 6102 474618 41546 475174
rect 42102 474618 77546 475174
rect 78102 474618 113546 475174
rect 114102 474618 149546 475174
rect 150102 474618 185546 475174
rect 186102 474618 221546 475174
rect 222102 474618 257546 475174
rect 258102 474618 293546 475174
rect 294102 474618 329546 475174
rect 330102 474618 365546 475174
rect 366102 474618 401546 475174
rect 402102 474618 437546 475174
rect 438102 474618 473546 475174
rect 474102 474618 509546 475174
rect 510102 474618 545546 475174
rect 546102 474618 581546 475174
rect 582102 474618 587262 475174
rect 587818 474618 588810 475174
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 470898 -1974 471454
rect -1418 470898 1826 471454
rect 2382 470898 37826 471454
rect 38382 470898 73826 471454
rect 74382 470898 109826 471454
rect 110382 470898 145826 471454
rect 146382 470898 181826 471454
rect 182382 470898 217826 471454
rect 218382 470898 253826 471454
rect 254382 470898 289826 471454
rect 290382 470898 325826 471454
rect 326382 470898 361826 471454
rect 362382 470898 397826 471454
rect 398382 470898 433826 471454
rect 434382 470898 469826 471454
rect 470382 470898 505826 471454
rect 506382 470898 541826 471454
rect 542382 470898 577826 471454
rect 578382 470898 585342 471454
rect 585898 470898 586890 471454
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464058 -8694 464614
rect -8138 464058 30986 464614
rect 31542 464058 66986 464614
rect 67542 464058 102986 464614
rect 103542 464058 138986 464614
rect 139542 464058 174986 464614
rect 175542 464058 210986 464614
rect 211542 464058 246986 464614
rect 247542 464058 282986 464614
rect 283542 464058 318986 464614
rect 319542 464058 354986 464614
rect 355542 464058 390986 464614
rect 391542 464058 426986 464614
rect 427542 464058 462986 464614
rect 463542 464058 498986 464614
rect 499542 464058 534986 464614
rect 535542 464058 570986 464614
rect 571542 464058 592062 464614
rect 592618 464058 592650 464614
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460338 -6774 460894
rect -6218 460338 27266 460894
rect 27822 460338 63266 460894
rect 63822 460338 99266 460894
rect 99822 460338 135266 460894
rect 135822 460338 171266 460894
rect 171822 460338 207266 460894
rect 207822 460338 243266 460894
rect 243822 460338 279266 460894
rect 279822 460338 315266 460894
rect 315822 460338 351266 460894
rect 351822 460338 387266 460894
rect 387822 460338 423266 460894
rect 423822 460338 459266 460894
rect 459822 460338 495266 460894
rect 495822 460338 531266 460894
rect 531822 460338 567266 460894
rect 567822 460338 590142 460894
rect 590698 460338 590730 460894
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456618 -4854 457174
rect -4298 456618 23546 457174
rect 24102 456618 59546 457174
rect 60102 456618 95546 457174
rect 96102 456618 131546 457174
rect 132102 456618 167546 457174
rect 168102 456618 203546 457174
rect 204102 456618 239546 457174
rect 240102 456618 275546 457174
rect 276102 456618 311546 457174
rect 312102 456618 347546 457174
rect 348102 456618 383546 457174
rect 384102 456618 419546 457174
rect 420102 456618 455546 457174
rect 456102 456618 491546 457174
rect 492102 456618 527546 457174
rect 528102 456618 563546 457174
rect 564102 456618 588222 457174
rect 588778 456618 588810 457174
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 452898 -2934 453454
rect -2378 452898 19826 453454
rect 20382 452898 55826 453454
rect 56382 452898 91826 453454
rect 92382 452898 127826 453454
rect 128382 452898 163826 453454
rect 164382 452898 199826 453454
rect 200382 452898 235826 453454
rect 236382 452898 271826 453454
rect 272382 452898 307826 453454
rect 308382 452898 343826 453454
rect 344382 452898 379826 453454
rect 380382 452898 415826 453454
rect 416382 452898 451826 453454
rect 452382 452898 487826 453454
rect 488382 452898 523826 453454
rect 524382 452898 559826 453454
rect 560382 452898 586302 453454
rect 586858 452898 586890 453454
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446058 -7734 446614
rect -7178 446058 12986 446614
rect 13542 446058 48986 446614
rect 49542 446058 84986 446614
rect 85542 446058 120986 446614
rect 121542 446058 156986 446614
rect 157542 446058 192986 446614
rect 193542 446058 228986 446614
rect 229542 446058 264986 446614
rect 265542 446058 300986 446614
rect 301542 446058 336986 446614
rect 337542 446058 372986 446614
rect 373542 446058 408986 446614
rect 409542 446058 444986 446614
rect 445542 446058 480986 446614
rect 481542 446058 516986 446614
rect 517542 446058 552986 446614
rect 553542 446058 591102 446614
rect 591658 446058 592650 446614
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442338 -5814 442894
rect -5258 442338 9266 442894
rect 9822 442338 45266 442894
rect 45822 442338 81266 442894
rect 81822 442338 117266 442894
rect 117822 442338 153266 442894
rect 153822 442338 189266 442894
rect 189822 442338 225266 442894
rect 225822 442338 261266 442894
rect 261822 442338 297266 442894
rect 297822 442338 333266 442894
rect 333822 442338 369266 442894
rect 369822 442338 405266 442894
rect 405822 442338 441266 442894
rect 441822 442338 477266 442894
rect 477822 442338 513266 442894
rect 513822 442338 549266 442894
rect 549822 442338 589182 442894
rect 589738 442338 590730 442894
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438618 -3894 439174
rect -3338 438618 5546 439174
rect 6102 438618 41546 439174
rect 42102 438618 77546 439174
rect 78102 438618 113546 439174
rect 114102 438618 149546 439174
rect 150102 438618 185546 439174
rect 186102 438618 221546 439174
rect 222102 438618 257546 439174
rect 258102 438618 293546 439174
rect 294102 438618 329546 439174
rect 330102 438618 365546 439174
rect 366102 438618 401546 439174
rect 402102 438618 437546 439174
rect 438102 438618 473546 439174
rect 474102 438618 509546 439174
rect 510102 438618 545546 439174
rect 546102 438618 581546 439174
rect 582102 438618 587262 439174
rect 587818 438618 588810 439174
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 434898 -1974 435454
rect -1418 434898 1826 435454
rect 2382 434898 37826 435454
rect 38382 434898 73826 435454
rect 74382 434898 109826 435454
rect 110382 434898 145826 435454
rect 146382 434898 181826 435454
rect 182382 434898 217826 435454
rect 218382 434898 253826 435454
rect 254382 434898 289826 435454
rect 290382 434898 325826 435454
rect 326382 434898 361826 435454
rect 362382 434898 397826 435454
rect 398382 434898 433826 435454
rect 434382 434898 469826 435454
rect 470382 434898 505826 435454
rect 506382 434898 541826 435454
rect 542382 434898 577826 435454
rect 578382 434898 585342 435454
rect 585898 434898 586890 435454
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428058 -8694 428614
rect -8138 428058 30986 428614
rect 31542 428058 66986 428614
rect 67542 428058 102986 428614
rect 103542 428058 138986 428614
rect 139542 428058 174986 428614
rect 175542 428058 210986 428614
rect 211542 428058 246986 428614
rect 247542 428058 282986 428614
rect 283542 428058 318986 428614
rect 319542 428058 354986 428614
rect 355542 428058 390986 428614
rect 391542 428058 426986 428614
rect 427542 428058 462986 428614
rect 463542 428058 498986 428614
rect 499542 428058 534986 428614
rect 535542 428058 570986 428614
rect 571542 428058 592062 428614
rect 592618 428058 592650 428614
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424338 -6774 424894
rect -6218 424338 27266 424894
rect 27822 424338 63266 424894
rect 63822 424338 99266 424894
rect 99822 424338 135266 424894
rect 135822 424338 171266 424894
rect 171822 424338 207266 424894
rect 207822 424338 243266 424894
rect 243822 424338 279266 424894
rect 279822 424338 315266 424894
rect 315822 424338 351266 424894
rect 351822 424338 387266 424894
rect 387822 424338 423266 424894
rect 423822 424338 459266 424894
rect 459822 424338 495266 424894
rect 495822 424338 531266 424894
rect 531822 424338 567266 424894
rect 567822 424338 590142 424894
rect 590698 424338 590730 424894
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420618 -4854 421174
rect -4298 420618 23546 421174
rect 24102 420618 59546 421174
rect 60102 420618 95546 421174
rect 96102 420618 131546 421174
rect 132102 420618 167546 421174
rect 168102 420618 203546 421174
rect 204102 420618 239546 421174
rect 240102 420618 275546 421174
rect 276102 420618 311546 421174
rect 312102 420618 347546 421174
rect 348102 420618 383546 421174
rect 384102 420618 419546 421174
rect 420102 420618 455546 421174
rect 456102 420618 491546 421174
rect 492102 420618 527546 421174
rect 528102 420618 563546 421174
rect 564102 420618 588222 421174
rect 588778 420618 588810 421174
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 416898 -2934 417454
rect -2378 416898 19826 417454
rect 20382 416898 55826 417454
rect 56382 416898 91826 417454
rect 92382 416898 127826 417454
rect 128382 416898 163826 417454
rect 164382 416898 199826 417454
rect 200382 416898 235826 417454
rect 236382 416898 271826 417454
rect 272382 416898 307826 417454
rect 308382 416898 343826 417454
rect 344382 416898 379826 417454
rect 380382 416898 415826 417454
rect 416382 416898 451826 417454
rect 452382 416898 487826 417454
rect 488382 416898 523826 417454
rect 524382 416898 559826 417454
rect 560382 416898 586302 417454
rect 586858 416898 586890 417454
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410058 -7734 410614
rect -7178 410058 12986 410614
rect 13542 410058 48986 410614
rect 49542 410058 84986 410614
rect 85542 410058 120986 410614
rect 121542 410058 156986 410614
rect 157542 410058 192986 410614
rect 193542 410058 228986 410614
rect 229542 410058 264986 410614
rect 265542 410058 300986 410614
rect 301542 410058 336986 410614
rect 337542 410058 372986 410614
rect 373542 410058 408986 410614
rect 409542 410058 444986 410614
rect 445542 410058 480986 410614
rect 481542 410058 516986 410614
rect 517542 410058 552986 410614
rect 553542 410058 591102 410614
rect 591658 410058 592650 410614
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406338 -5814 406894
rect -5258 406338 9266 406894
rect 9822 406338 45266 406894
rect 45822 406338 81266 406894
rect 81822 406338 117266 406894
rect 117822 406338 153266 406894
rect 153822 406338 189266 406894
rect 189822 406338 225266 406894
rect 225822 406338 261266 406894
rect 261822 406338 297266 406894
rect 297822 406338 333266 406894
rect 333822 406338 369266 406894
rect 369822 406338 405266 406894
rect 405822 406338 441266 406894
rect 441822 406338 477266 406894
rect 477822 406338 513266 406894
rect 513822 406338 549266 406894
rect 549822 406338 589182 406894
rect 589738 406338 590730 406894
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402618 -3894 403174
rect -3338 402618 5546 403174
rect 6102 402618 41546 403174
rect 42102 402618 77546 403174
rect 78102 402618 113546 403174
rect 114102 402618 149546 403174
rect 150102 402618 185546 403174
rect 186102 402618 221546 403174
rect 222102 402618 257546 403174
rect 258102 402618 293546 403174
rect 294102 402618 329546 403174
rect 330102 402618 365546 403174
rect 366102 402618 401546 403174
rect 402102 402618 437546 403174
rect 438102 402618 473546 403174
rect 474102 402618 509546 403174
rect 510102 402618 545546 403174
rect 546102 402618 581546 403174
rect 582102 402618 587262 403174
rect 587818 402618 588810 403174
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 398898 -1974 399454
rect -1418 398898 1826 399454
rect 2382 398898 37826 399454
rect 38382 398898 73826 399454
rect 74382 398898 109826 399454
rect 110382 398898 145826 399454
rect 146382 398898 181826 399454
rect 182382 398898 217826 399454
rect 218382 398898 253826 399454
rect 254382 398898 289826 399454
rect 290382 398898 325826 399454
rect 326382 398898 361826 399454
rect 362382 398898 397826 399454
rect 398382 398898 433826 399454
rect 434382 398898 469826 399454
rect 470382 398898 505826 399454
rect 506382 398898 541826 399454
rect 542382 398898 577826 399454
rect 578382 398898 585342 399454
rect 585898 398898 586890 399454
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392058 -8694 392614
rect -8138 392058 30986 392614
rect 31542 392058 66986 392614
rect 67542 392058 102986 392614
rect 103542 392058 138986 392614
rect 139542 392058 174986 392614
rect 175542 392058 210986 392614
rect 211542 392058 246986 392614
rect 247542 392058 282986 392614
rect 283542 392058 318986 392614
rect 319542 392058 354986 392614
rect 355542 392058 390986 392614
rect 391542 392058 426986 392614
rect 427542 392058 462986 392614
rect 463542 392058 498986 392614
rect 499542 392058 534986 392614
rect 535542 392058 570986 392614
rect 571542 392058 592062 392614
rect 592618 392058 592650 392614
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388338 -6774 388894
rect -6218 388338 27266 388894
rect 27822 388338 63266 388894
rect 63822 388338 99266 388894
rect 99822 388338 135266 388894
rect 135822 388338 171266 388894
rect 171822 388338 207266 388894
rect 207822 388338 243266 388894
rect 243822 388338 279266 388894
rect 279822 388338 315266 388894
rect 315822 388338 351266 388894
rect 351822 388338 387266 388894
rect 387822 388338 423266 388894
rect 423822 388338 459266 388894
rect 459822 388338 495266 388894
rect 495822 388338 531266 388894
rect 531822 388338 567266 388894
rect 567822 388338 590142 388894
rect 590698 388338 590730 388894
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384618 -4854 385174
rect -4298 384618 23546 385174
rect 24102 384618 59546 385174
rect 60102 384618 95546 385174
rect 96102 384618 131546 385174
rect 132102 384618 167546 385174
rect 168102 384618 203546 385174
rect 204102 384618 239546 385174
rect 240102 384618 275546 385174
rect 276102 384618 311546 385174
rect 312102 384618 347546 385174
rect 348102 384618 383546 385174
rect 384102 384618 419546 385174
rect 420102 384618 455546 385174
rect 456102 384618 491546 385174
rect 492102 384618 527546 385174
rect 528102 384618 563546 385174
rect 564102 384618 588222 385174
rect 588778 384618 588810 385174
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 380898 -2934 381454
rect -2378 380898 19826 381454
rect 20382 380898 55826 381454
rect 56382 380898 91826 381454
rect 92382 380898 127826 381454
rect 128382 380898 163826 381454
rect 164382 380898 199826 381454
rect 200382 380898 235826 381454
rect 236382 380898 271826 381454
rect 272382 380898 307826 381454
rect 308382 380898 343826 381454
rect 344382 380898 379826 381454
rect 380382 380898 415826 381454
rect 416382 380898 451826 381454
rect 452382 380898 487826 381454
rect 488382 380898 523826 381454
rect 524382 380898 559826 381454
rect 560382 380898 586302 381454
rect 586858 380898 586890 381454
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374058 -7734 374614
rect -7178 374058 12986 374614
rect 13542 374058 48986 374614
rect 49542 374058 84986 374614
rect 85542 374058 120986 374614
rect 121542 374058 156986 374614
rect 157542 374058 192986 374614
rect 193542 374058 228986 374614
rect 229542 374058 300986 374614
rect 301542 374058 336986 374614
rect 337542 374058 372986 374614
rect 373542 374058 408986 374614
rect 409542 374058 444986 374614
rect 445542 374058 480986 374614
rect 481542 374058 516986 374614
rect 517542 374058 552986 374614
rect 553542 374058 591102 374614
rect 591658 374058 592650 374614
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370338 -5814 370894
rect -5258 370338 9266 370894
rect 9822 370338 45266 370894
rect 45822 370338 81266 370894
rect 81822 370338 117266 370894
rect 117822 370338 153266 370894
rect 153822 370338 189266 370894
rect 189822 370338 225266 370894
rect 225822 370338 297266 370894
rect 297822 370338 333266 370894
rect 333822 370338 369266 370894
rect 369822 370338 405266 370894
rect 405822 370338 441266 370894
rect 441822 370338 477266 370894
rect 477822 370338 513266 370894
rect 513822 370338 549266 370894
rect 549822 370338 589182 370894
rect 589738 370338 590730 370894
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366618 -3894 367174
rect -3338 366618 5546 367174
rect 6102 366618 41546 367174
rect 42102 366618 77546 367174
rect 78102 366618 113546 367174
rect 114102 366618 149546 367174
rect 150102 366618 185546 367174
rect 186102 366618 221546 367174
rect 222102 366618 329546 367174
rect 330102 366618 365546 367174
rect 366102 366618 401546 367174
rect 402102 366618 437546 367174
rect 438102 366618 473546 367174
rect 474102 366618 509546 367174
rect 510102 366618 545546 367174
rect 546102 366618 581546 367174
rect 582102 366618 587262 367174
rect 587818 366618 588810 367174
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 362898 -1974 363454
rect -1418 362898 1826 363454
rect 2382 362898 37826 363454
rect 38382 362898 73826 363454
rect 74382 362898 109826 363454
rect 110382 362898 145826 363454
rect 146382 362898 181826 363454
rect 182382 362898 217826 363454
rect 218382 363218 239250 363454
rect 239486 363218 269970 363454
rect 270206 363218 325826 363454
rect 218382 363134 325826 363218
rect 218382 362898 239250 363134
rect 239486 362898 269970 363134
rect 270206 362898 325826 363134
rect 326382 362898 361826 363454
rect 362382 362898 397826 363454
rect 398382 362898 433826 363454
rect 434382 362898 469826 363454
rect 470382 362898 505826 363454
rect 506382 362898 541826 363454
rect 542382 362898 577826 363454
rect 578382 362898 585342 363454
rect 585898 362898 586890 363454
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356058 -8694 356614
rect -8138 356058 30986 356614
rect 31542 356058 66986 356614
rect 67542 356058 102986 356614
rect 103542 356058 138986 356614
rect 139542 356058 174986 356614
rect 175542 356058 210986 356614
rect 211542 356058 318986 356614
rect 319542 356058 354986 356614
rect 355542 356058 390986 356614
rect 391542 356058 426986 356614
rect 427542 356058 462986 356614
rect 463542 356058 498986 356614
rect 499542 356058 534986 356614
rect 535542 356058 570986 356614
rect 571542 356058 592062 356614
rect 592618 356058 592650 356614
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352338 -6774 352894
rect -6218 352338 27266 352894
rect 27822 352338 63266 352894
rect 63822 352338 99266 352894
rect 99822 352338 135266 352894
rect 135822 352338 171266 352894
rect 171822 352338 207266 352894
rect 207822 352338 315266 352894
rect 315822 352338 351266 352894
rect 351822 352338 387266 352894
rect 387822 352338 423266 352894
rect 423822 352338 459266 352894
rect 459822 352338 495266 352894
rect 495822 352338 531266 352894
rect 531822 352338 567266 352894
rect 567822 352338 590142 352894
rect 590698 352338 590730 352894
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348618 -4854 349174
rect -4298 348618 23546 349174
rect 24102 348618 59546 349174
rect 60102 348618 95546 349174
rect 96102 348618 131546 349174
rect 132102 348618 167546 349174
rect 168102 348618 203546 349174
rect 204102 348618 311546 349174
rect 312102 348618 347546 349174
rect 348102 348618 383546 349174
rect 384102 348618 419546 349174
rect 420102 348618 455546 349174
rect 456102 348618 491546 349174
rect 492102 348618 527546 349174
rect 528102 348618 563546 349174
rect 564102 348618 588222 349174
rect 588778 348618 588810 349174
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 344898 -2934 345454
rect -2378 344898 19826 345454
rect 20382 344898 55826 345454
rect 56382 344898 91826 345454
rect 92382 344898 127826 345454
rect 128382 344898 163826 345454
rect 164382 344898 199826 345454
rect 200382 345218 254610 345454
rect 254846 345218 285330 345454
rect 285566 345218 307826 345454
rect 200382 345134 307826 345218
rect 200382 344898 254610 345134
rect 254846 344898 285330 345134
rect 285566 344898 307826 345134
rect 308382 344898 343826 345454
rect 344382 344898 379826 345454
rect 380382 344898 415826 345454
rect 416382 344898 451826 345454
rect 452382 344898 487826 345454
rect 488382 344898 523826 345454
rect 524382 344898 559826 345454
rect 560382 344898 586302 345454
rect 586858 344898 586890 345454
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338058 -7734 338614
rect -7178 338058 12986 338614
rect 13542 338058 48986 338614
rect 49542 338058 84986 338614
rect 85542 338058 120986 338614
rect 121542 338058 156986 338614
rect 157542 338058 192986 338614
rect 193542 338058 228986 338614
rect 229542 338058 300986 338614
rect 301542 338058 336986 338614
rect 337542 338058 372986 338614
rect 373542 338058 408986 338614
rect 409542 338058 444986 338614
rect 445542 338058 480986 338614
rect 481542 338058 516986 338614
rect 517542 338058 552986 338614
rect 553542 338058 591102 338614
rect 591658 338058 592650 338614
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334338 -5814 334894
rect -5258 334338 9266 334894
rect 9822 334338 45266 334894
rect 45822 334338 81266 334894
rect 81822 334338 117266 334894
rect 117822 334338 153266 334894
rect 153822 334338 189266 334894
rect 189822 334338 225266 334894
rect 225822 334338 261266 334894
rect 261822 334338 297266 334894
rect 297822 334338 333266 334894
rect 333822 334338 369266 334894
rect 369822 334338 405266 334894
rect 405822 334338 441266 334894
rect 441822 334338 477266 334894
rect 477822 334338 513266 334894
rect 513822 334338 549266 334894
rect 549822 334338 589182 334894
rect 589738 334338 590730 334894
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330618 -3894 331174
rect -3338 330618 5546 331174
rect 6102 330618 41546 331174
rect 42102 330618 77546 331174
rect 78102 330618 113546 331174
rect 114102 330618 149546 331174
rect 150102 330618 185546 331174
rect 186102 330618 221546 331174
rect 222102 330618 257546 331174
rect 258102 330618 293546 331174
rect 294102 330618 329546 331174
rect 330102 330618 365546 331174
rect 366102 330618 401546 331174
rect 402102 330618 437546 331174
rect 438102 330618 473546 331174
rect 474102 330618 509546 331174
rect 510102 330618 545546 331174
rect 546102 330618 581546 331174
rect 582102 330618 587262 331174
rect 587818 330618 588810 331174
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 326898 -1974 327454
rect -1418 326898 1826 327454
rect 2382 326898 37826 327454
rect 38382 326898 73826 327454
rect 74382 326898 109826 327454
rect 110382 326898 145826 327454
rect 146382 326898 181826 327454
rect 182382 326898 217826 327454
rect 218382 326898 253826 327454
rect 254382 326898 289826 327454
rect 290382 326898 325826 327454
rect 326382 326898 361826 327454
rect 362382 326898 397826 327454
rect 398382 326898 433826 327454
rect 434382 326898 469826 327454
rect 470382 326898 505826 327454
rect 506382 326898 541826 327454
rect 542382 326898 577826 327454
rect 578382 326898 585342 327454
rect 585898 326898 586890 327454
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320058 -8694 320614
rect -8138 320058 30986 320614
rect 31542 320058 66986 320614
rect 67542 320058 102986 320614
rect 103542 320058 138986 320614
rect 139542 320058 174986 320614
rect 175542 320058 210986 320614
rect 211542 320058 246986 320614
rect 247542 320058 282986 320614
rect 283542 320058 318986 320614
rect 319542 320058 354986 320614
rect 355542 320058 390986 320614
rect 391542 320058 426986 320614
rect 427542 320058 462986 320614
rect 463542 320058 498986 320614
rect 499542 320058 534986 320614
rect 535542 320058 570986 320614
rect 571542 320058 592062 320614
rect 592618 320058 592650 320614
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316338 -6774 316894
rect -6218 316338 27266 316894
rect 27822 316338 63266 316894
rect 63822 316338 99266 316894
rect 99822 316338 135266 316894
rect 135822 316338 171266 316894
rect 171822 316338 207266 316894
rect 207822 316338 243266 316894
rect 243822 316338 279266 316894
rect 279822 316338 315266 316894
rect 315822 316338 351266 316894
rect 351822 316338 387266 316894
rect 387822 316338 423266 316894
rect 423822 316338 459266 316894
rect 459822 316338 495266 316894
rect 495822 316338 531266 316894
rect 531822 316338 567266 316894
rect 567822 316338 590142 316894
rect 590698 316338 590730 316894
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312618 -4854 313174
rect -4298 312618 23546 313174
rect 24102 312618 59546 313174
rect 60102 312618 95546 313174
rect 96102 312618 131546 313174
rect 132102 312618 167546 313174
rect 168102 312618 203546 313174
rect 204102 312618 239546 313174
rect 240102 312618 275546 313174
rect 276102 312618 311546 313174
rect 312102 312618 347546 313174
rect 348102 312618 383546 313174
rect 384102 312618 419546 313174
rect 420102 312618 455546 313174
rect 456102 312618 491546 313174
rect 492102 312618 527546 313174
rect 528102 312618 563546 313174
rect 564102 312618 588222 313174
rect 588778 312618 588810 313174
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 308898 -2934 309454
rect -2378 308898 19826 309454
rect 20382 308898 55826 309454
rect 56382 308898 91826 309454
rect 92382 308898 127826 309454
rect 128382 308898 163826 309454
rect 164382 308898 199826 309454
rect 200382 308898 235826 309454
rect 236382 308898 271826 309454
rect 272382 308898 307826 309454
rect 308382 308898 343826 309454
rect 344382 308898 379826 309454
rect 380382 308898 415826 309454
rect 416382 308898 451826 309454
rect 452382 308898 487826 309454
rect 488382 308898 523826 309454
rect 524382 308898 559826 309454
rect 560382 308898 586302 309454
rect 586858 308898 586890 309454
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302058 -7734 302614
rect -7178 302058 12986 302614
rect 13542 302058 48986 302614
rect 49542 302058 84986 302614
rect 85542 302058 120986 302614
rect 121542 302058 156986 302614
rect 157542 302058 192986 302614
rect 193542 302058 228986 302614
rect 229542 302058 264986 302614
rect 265542 302058 300986 302614
rect 301542 302058 336986 302614
rect 337542 302058 372986 302614
rect 373542 302058 408986 302614
rect 409542 302058 444986 302614
rect 445542 302058 480986 302614
rect 481542 302058 516986 302614
rect 517542 302058 552986 302614
rect 553542 302058 591102 302614
rect 591658 302058 592650 302614
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298338 -5814 298894
rect -5258 298338 9266 298894
rect 9822 298338 45266 298894
rect 45822 298338 81266 298894
rect 81822 298338 117266 298894
rect 117822 298338 153266 298894
rect 153822 298338 189266 298894
rect 189822 298338 225266 298894
rect 225822 298338 261266 298894
rect 261822 298338 297266 298894
rect 297822 298338 333266 298894
rect 333822 298338 369266 298894
rect 369822 298338 405266 298894
rect 405822 298338 441266 298894
rect 441822 298338 477266 298894
rect 477822 298338 513266 298894
rect 513822 298338 549266 298894
rect 549822 298338 589182 298894
rect 589738 298338 590730 298894
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294618 -3894 295174
rect -3338 294618 5546 295174
rect 6102 294618 41546 295174
rect 42102 294618 77546 295174
rect 78102 294618 113546 295174
rect 114102 294618 149546 295174
rect 150102 294618 185546 295174
rect 186102 294618 221546 295174
rect 222102 294618 257546 295174
rect 258102 294618 293546 295174
rect 294102 294618 329546 295174
rect 330102 294618 365546 295174
rect 366102 294618 401546 295174
rect 402102 294618 437546 295174
rect 438102 294618 473546 295174
rect 474102 294618 509546 295174
rect 510102 294618 545546 295174
rect 546102 294618 581546 295174
rect 582102 294618 587262 295174
rect 587818 294618 588810 295174
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 290898 -1974 291454
rect -1418 290898 1826 291454
rect 2382 290898 37826 291454
rect 38382 290898 73826 291454
rect 74382 290898 109826 291454
rect 110382 290898 145826 291454
rect 146382 290898 181826 291454
rect 182382 290898 217826 291454
rect 218382 290898 253826 291454
rect 254382 290898 289826 291454
rect 290382 290898 325826 291454
rect 326382 290898 361826 291454
rect 362382 290898 397826 291454
rect 398382 290898 433826 291454
rect 434382 290898 469826 291454
rect 470382 290898 505826 291454
rect 506382 290898 541826 291454
rect 542382 290898 577826 291454
rect 578382 290898 585342 291454
rect 585898 290898 586890 291454
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284058 -8694 284614
rect -8138 284058 30986 284614
rect 31542 284058 66986 284614
rect 67542 284058 102986 284614
rect 103542 284058 138986 284614
rect 139542 284058 174986 284614
rect 175542 284058 210986 284614
rect 211542 284058 246986 284614
rect 247542 284058 282986 284614
rect 283542 284058 318986 284614
rect 319542 284058 354986 284614
rect 355542 284058 390986 284614
rect 391542 284058 426986 284614
rect 427542 284058 462986 284614
rect 463542 284058 498986 284614
rect 499542 284058 534986 284614
rect 535542 284058 570986 284614
rect 571542 284058 592062 284614
rect 592618 284058 592650 284614
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280338 -6774 280894
rect -6218 280338 27266 280894
rect 27822 280338 63266 280894
rect 63822 280338 99266 280894
rect 99822 280338 135266 280894
rect 135822 280338 171266 280894
rect 171822 280338 207266 280894
rect 207822 280338 243266 280894
rect 243822 280338 279266 280894
rect 279822 280338 315266 280894
rect 315822 280338 351266 280894
rect 351822 280338 387266 280894
rect 387822 280338 423266 280894
rect 423822 280338 459266 280894
rect 459822 280338 495266 280894
rect 495822 280338 531266 280894
rect 531822 280338 567266 280894
rect 567822 280338 590142 280894
rect 590698 280338 590730 280894
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276618 -4854 277174
rect -4298 276618 23546 277174
rect 24102 276618 59546 277174
rect 60102 276618 95546 277174
rect 96102 276618 131546 277174
rect 132102 276618 167546 277174
rect 168102 276618 203546 277174
rect 204102 276618 239546 277174
rect 240102 276618 275546 277174
rect 276102 276618 311546 277174
rect 312102 276618 347546 277174
rect 348102 276618 383546 277174
rect 384102 276618 419546 277174
rect 420102 276618 455546 277174
rect 456102 276618 491546 277174
rect 492102 276618 527546 277174
rect 528102 276618 563546 277174
rect 564102 276618 588222 277174
rect 588778 276618 588810 277174
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 272898 -2934 273454
rect -2378 272898 19826 273454
rect 20382 272898 55826 273454
rect 56382 272898 91826 273454
rect 92382 272898 127826 273454
rect 128382 272898 163826 273454
rect 164382 272898 199826 273454
rect 200382 272898 235826 273454
rect 236382 272898 271826 273454
rect 272382 272898 307826 273454
rect 308382 272898 343826 273454
rect 344382 272898 379826 273454
rect 380382 272898 415826 273454
rect 416382 272898 451826 273454
rect 452382 272898 487826 273454
rect 488382 272898 523826 273454
rect 524382 272898 559826 273454
rect 560382 272898 586302 273454
rect 586858 272898 586890 273454
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266058 -7734 266614
rect -7178 266058 12986 266614
rect 13542 266058 48986 266614
rect 49542 266058 84986 266614
rect 85542 266058 120986 266614
rect 121542 266058 156986 266614
rect 157542 266058 192986 266614
rect 193542 266058 228986 266614
rect 229542 266058 264986 266614
rect 265542 266058 300986 266614
rect 301542 266058 336986 266614
rect 337542 266058 372986 266614
rect 373542 266058 408986 266614
rect 409542 266058 444986 266614
rect 445542 266058 480986 266614
rect 481542 266058 516986 266614
rect 517542 266058 552986 266614
rect 553542 266058 591102 266614
rect 591658 266058 592650 266614
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262338 -5814 262894
rect -5258 262338 9266 262894
rect 9822 262338 45266 262894
rect 45822 262338 81266 262894
rect 81822 262338 117266 262894
rect 117822 262338 153266 262894
rect 153822 262338 189266 262894
rect 189822 262338 225266 262894
rect 225822 262338 261266 262894
rect 261822 262338 297266 262894
rect 297822 262338 333266 262894
rect 333822 262338 369266 262894
rect 369822 262338 405266 262894
rect 405822 262338 441266 262894
rect 441822 262338 477266 262894
rect 477822 262338 513266 262894
rect 513822 262338 549266 262894
rect 549822 262338 589182 262894
rect 589738 262338 590730 262894
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258618 -3894 259174
rect -3338 258618 5546 259174
rect 6102 258618 41546 259174
rect 42102 258618 77546 259174
rect 78102 258618 113546 259174
rect 114102 258618 149546 259174
rect 150102 258618 185546 259174
rect 186102 258618 221546 259174
rect 222102 258618 257546 259174
rect 258102 258618 293546 259174
rect 294102 258618 329546 259174
rect 330102 258618 365546 259174
rect 366102 258618 401546 259174
rect 402102 258618 437546 259174
rect 438102 258618 473546 259174
rect 474102 258618 509546 259174
rect 510102 258618 545546 259174
rect 546102 258618 581546 259174
rect 582102 258618 587262 259174
rect 587818 258618 588810 259174
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 254898 -1974 255454
rect -1418 254898 1826 255454
rect 2382 254898 37826 255454
rect 38382 254898 73826 255454
rect 74382 254898 109826 255454
rect 110382 254898 145826 255454
rect 146382 254898 181826 255454
rect 182382 254898 217826 255454
rect 218382 254898 253826 255454
rect 254382 254898 289826 255454
rect 290382 254898 325826 255454
rect 326382 254898 361826 255454
rect 362382 254898 397826 255454
rect 398382 254898 433826 255454
rect 434382 254898 469826 255454
rect 470382 254898 505826 255454
rect 506382 254898 541826 255454
rect 542382 254898 577826 255454
rect 578382 254898 585342 255454
rect 585898 254898 586890 255454
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248058 -8694 248614
rect -8138 248058 30986 248614
rect 31542 248058 66986 248614
rect 67542 248058 102986 248614
rect 103542 248058 138986 248614
rect 139542 248058 174986 248614
rect 175542 248058 210986 248614
rect 211542 248058 246986 248614
rect 247542 248058 282986 248614
rect 283542 248058 318986 248614
rect 319542 248058 354986 248614
rect 355542 248058 390986 248614
rect 391542 248058 426986 248614
rect 427542 248058 462986 248614
rect 463542 248058 498986 248614
rect 499542 248058 534986 248614
rect 535542 248058 570986 248614
rect 571542 248058 592062 248614
rect 592618 248058 592650 248614
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244338 -6774 244894
rect -6218 244338 27266 244894
rect 27822 244338 63266 244894
rect 63822 244338 99266 244894
rect 99822 244338 135266 244894
rect 135822 244338 171266 244894
rect 171822 244338 207266 244894
rect 207822 244338 243266 244894
rect 243822 244338 279266 244894
rect 279822 244338 315266 244894
rect 315822 244338 351266 244894
rect 351822 244338 387266 244894
rect 387822 244338 423266 244894
rect 423822 244338 459266 244894
rect 459822 244338 495266 244894
rect 495822 244338 531266 244894
rect 531822 244338 567266 244894
rect 567822 244338 590142 244894
rect 590698 244338 590730 244894
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240618 -4854 241174
rect -4298 240618 23546 241174
rect 24102 240618 59546 241174
rect 60102 240618 95546 241174
rect 96102 240618 131546 241174
rect 132102 240618 167546 241174
rect 168102 240618 203546 241174
rect 204102 240618 239546 241174
rect 240102 240618 275546 241174
rect 276102 240618 311546 241174
rect 312102 240618 347546 241174
rect 348102 240618 383546 241174
rect 384102 240618 419546 241174
rect 420102 240618 455546 241174
rect 456102 240618 491546 241174
rect 492102 240618 527546 241174
rect 528102 240618 563546 241174
rect 564102 240618 588222 241174
rect 588778 240618 588810 241174
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 236898 -2934 237454
rect -2378 236898 19826 237454
rect 20382 236898 55826 237454
rect 56382 236898 91826 237454
rect 92382 236898 127826 237454
rect 128382 236898 163826 237454
rect 164382 236898 199826 237454
rect 200382 236898 235826 237454
rect 236382 236898 271826 237454
rect 272382 236898 307826 237454
rect 308382 236898 343826 237454
rect 344382 236898 379826 237454
rect 380382 236898 415826 237454
rect 416382 236898 451826 237454
rect 452382 236898 487826 237454
rect 488382 236898 523826 237454
rect 524382 236898 559826 237454
rect 560382 236898 586302 237454
rect 586858 236898 586890 237454
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230058 -7734 230614
rect -7178 230058 12986 230614
rect 13542 230058 48986 230614
rect 49542 230058 84986 230614
rect 85542 230058 120986 230614
rect 121542 230058 156986 230614
rect 157542 230058 192986 230614
rect 193542 230058 228986 230614
rect 229542 230058 264986 230614
rect 265542 230058 300986 230614
rect 301542 230058 336986 230614
rect 337542 230058 372986 230614
rect 373542 230058 408986 230614
rect 409542 230058 444986 230614
rect 445542 230058 480986 230614
rect 481542 230058 516986 230614
rect 517542 230058 552986 230614
rect 553542 230058 591102 230614
rect 591658 230058 592650 230614
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226338 -5814 226894
rect -5258 226338 9266 226894
rect 9822 226338 45266 226894
rect 45822 226338 81266 226894
rect 81822 226338 117266 226894
rect 117822 226338 153266 226894
rect 153822 226338 189266 226894
rect 189822 226338 225266 226894
rect 225822 226338 261266 226894
rect 261822 226338 297266 226894
rect 297822 226338 333266 226894
rect 333822 226338 369266 226894
rect 369822 226338 405266 226894
rect 405822 226338 441266 226894
rect 441822 226338 477266 226894
rect 477822 226338 513266 226894
rect 513822 226338 549266 226894
rect 549822 226338 589182 226894
rect 589738 226338 590730 226894
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222618 -3894 223174
rect -3338 222618 5546 223174
rect 6102 222618 41546 223174
rect 42102 222618 77546 223174
rect 78102 222618 113546 223174
rect 114102 222618 149546 223174
rect 150102 222618 185546 223174
rect 186102 222618 221546 223174
rect 222102 222618 257546 223174
rect 258102 222618 293546 223174
rect 294102 222618 329546 223174
rect 330102 222618 365546 223174
rect 366102 222618 401546 223174
rect 402102 222618 437546 223174
rect 438102 222618 473546 223174
rect 474102 222618 509546 223174
rect 510102 222618 545546 223174
rect 546102 222618 581546 223174
rect 582102 222618 587262 223174
rect 587818 222618 588810 223174
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 218898 -1974 219454
rect -1418 218898 1826 219454
rect 2382 218898 37826 219454
rect 38382 218898 73826 219454
rect 74382 218898 109826 219454
rect 110382 218898 145826 219454
rect 146382 218898 181826 219454
rect 182382 218898 217826 219454
rect 218382 218898 253826 219454
rect 254382 218898 289826 219454
rect 290382 218898 325826 219454
rect 326382 218898 361826 219454
rect 362382 218898 397826 219454
rect 398382 218898 433826 219454
rect 434382 218898 469826 219454
rect 470382 218898 505826 219454
rect 506382 218898 541826 219454
rect 542382 218898 577826 219454
rect 578382 218898 585342 219454
rect 585898 218898 586890 219454
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212058 -8694 212614
rect -8138 212058 30986 212614
rect 31542 212058 66986 212614
rect 67542 212058 102986 212614
rect 103542 212058 138986 212614
rect 139542 212058 174986 212614
rect 175542 212058 210986 212614
rect 211542 212058 246986 212614
rect 247542 212058 282986 212614
rect 283542 212058 318986 212614
rect 319542 212058 354986 212614
rect 355542 212058 390986 212614
rect 391542 212058 426986 212614
rect 427542 212058 462986 212614
rect 463542 212058 498986 212614
rect 499542 212058 534986 212614
rect 535542 212058 570986 212614
rect 571542 212058 592062 212614
rect 592618 212058 592650 212614
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208338 -6774 208894
rect -6218 208338 27266 208894
rect 27822 208338 63266 208894
rect 63822 208338 99266 208894
rect 99822 208338 135266 208894
rect 135822 208338 171266 208894
rect 171822 208338 207266 208894
rect 207822 208338 243266 208894
rect 243822 208338 279266 208894
rect 279822 208338 315266 208894
rect 315822 208338 351266 208894
rect 351822 208338 387266 208894
rect 387822 208338 423266 208894
rect 423822 208338 459266 208894
rect 459822 208338 495266 208894
rect 495822 208338 531266 208894
rect 531822 208338 567266 208894
rect 567822 208338 590142 208894
rect 590698 208338 590730 208894
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204618 -4854 205174
rect -4298 204618 23546 205174
rect 24102 204618 59546 205174
rect 60102 204618 95546 205174
rect 96102 204618 131546 205174
rect 132102 204618 167546 205174
rect 168102 204618 203546 205174
rect 204102 204618 239546 205174
rect 240102 204618 275546 205174
rect 276102 204618 311546 205174
rect 312102 204618 347546 205174
rect 348102 204618 383546 205174
rect 384102 204618 419546 205174
rect 420102 204618 455546 205174
rect 456102 204618 491546 205174
rect 492102 204618 527546 205174
rect 528102 204618 563546 205174
rect 564102 204618 588222 205174
rect 588778 204618 588810 205174
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 200898 -2934 201454
rect -2378 200898 19826 201454
rect 20382 200898 55826 201454
rect 56382 200898 91826 201454
rect 92382 200898 127826 201454
rect 128382 200898 163826 201454
rect 164382 200898 199826 201454
rect 200382 200898 235826 201454
rect 236382 200898 271826 201454
rect 272382 200898 307826 201454
rect 308382 200898 343826 201454
rect 344382 200898 379826 201454
rect 380382 200898 415826 201454
rect 416382 200898 451826 201454
rect 452382 200898 487826 201454
rect 488382 200898 523826 201454
rect 524382 200898 559826 201454
rect 560382 200898 586302 201454
rect 586858 200898 586890 201454
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194058 -7734 194614
rect -7178 194058 12986 194614
rect 13542 194058 48986 194614
rect 49542 194058 84986 194614
rect 85542 194058 120986 194614
rect 121542 194058 156986 194614
rect 157542 194058 192986 194614
rect 193542 194058 228986 194614
rect 229542 194058 264986 194614
rect 265542 194058 300986 194614
rect 301542 194058 336986 194614
rect 337542 194058 372986 194614
rect 373542 194058 408986 194614
rect 409542 194058 444986 194614
rect 445542 194058 480986 194614
rect 481542 194058 516986 194614
rect 517542 194058 552986 194614
rect 553542 194058 591102 194614
rect 591658 194058 592650 194614
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190338 -5814 190894
rect -5258 190338 9266 190894
rect 9822 190338 45266 190894
rect 45822 190338 81266 190894
rect 81822 190338 117266 190894
rect 117822 190338 153266 190894
rect 153822 190338 189266 190894
rect 189822 190338 225266 190894
rect 225822 190338 261266 190894
rect 261822 190338 297266 190894
rect 297822 190338 333266 190894
rect 333822 190338 369266 190894
rect 369822 190338 405266 190894
rect 405822 190338 441266 190894
rect 441822 190338 477266 190894
rect 477822 190338 513266 190894
rect 513822 190338 549266 190894
rect 549822 190338 589182 190894
rect 589738 190338 590730 190894
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186618 -3894 187174
rect -3338 186618 5546 187174
rect 6102 186618 41546 187174
rect 42102 186618 77546 187174
rect 78102 186618 113546 187174
rect 114102 186618 149546 187174
rect 150102 186618 185546 187174
rect 186102 186618 221546 187174
rect 222102 186618 257546 187174
rect 258102 186618 293546 187174
rect 294102 186618 329546 187174
rect 330102 186618 365546 187174
rect 366102 186618 401546 187174
rect 402102 186618 437546 187174
rect 438102 186618 473546 187174
rect 474102 186618 509546 187174
rect 510102 186618 545546 187174
rect 546102 186618 581546 187174
rect 582102 186618 587262 187174
rect 587818 186618 588810 187174
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 182898 -1974 183454
rect -1418 182898 1826 183454
rect 2382 182898 37826 183454
rect 38382 182898 73826 183454
rect 74382 182898 109826 183454
rect 110382 182898 145826 183454
rect 146382 182898 181826 183454
rect 182382 182898 217826 183454
rect 218382 182898 253826 183454
rect 254382 182898 289826 183454
rect 290382 182898 325826 183454
rect 326382 182898 361826 183454
rect 362382 182898 397826 183454
rect 398382 182898 433826 183454
rect 434382 182898 469826 183454
rect 470382 182898 505826 183454
rect 506382 182898 541826 183454
rect 542382 182898 577826 183454
rect 578382 182898 585342 183454
rect 585898 182898 586890 183454
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176058 -8694 176614
rect -8138 176058 30986 176614
rect 31542 176058 66986 176614
rect 67542 176058 102986 176614
rect 103542 176058 138986 176614
rect 139542 176058 174986 176614
rect 175542 176058 210986 176614
rect 211542 176058 246986 176614
rect 247542 176058 282986 176614
rect 283542 176058 318986 176614
rect 319542 176058 354986 176614
rect 355542 176058 390986 176614
rect 391542 176058 426986 176614
rect 427542 176058 462986 176614
rect 463542 176058 498986 176614
rect 499542 176058 534986 176614
rect 535542 176058 570986 176614
rect 571542 176058 592062 176614
rect 592618 176058 592650 176614
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172338 -6774 172894
rect -6218 172338 27266 172894
rect 27822 172338 63266 172894
rect 63822 172338 99266 172894
rect 99822 172338 135266 172894
rect 135822 172338 171266 172894
rect 171822 172338 207266 172894
rect 207822 172338 243266 172894
rect 243822 172338 279266 172894
rect 279822 172338 315266 172894
rect 315822 172338 351266 172894
rect 351822 172338 387266 172894
rect 387822 172338 423266 172894
rect 423822 172338 459266 172894
rect 459822 172338 495266 172894
rect 495822 172338 531266 172894
rect 531822 172338 567266 172894
rect 567822 172338 590142 172894
rect 590698 172338 590730 172894
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168618 -4854 169174
rect -4298 168618 23546 169174
rect 24102 168618 59546 169174
rect 60102 168618 95546 169174
rect 96102 168618 131546 169174
rect 132102 168618 167546 169174
rect 168102 168618 203546 169174
rect 204102 168618 239546 169174
rect 240102 168618 275546 169174
rect 276102 168618 311546 169174
rect 312102 168618 347546 169174
rect 348102 168618 383546 169174
rect 384102 168618 419546 169174
rect 420102 168618 455546 169174
rect 456102 168618 491546 169174
rect 492102 168618 527546 169174
rect 528102 168618 563546 169174
rect 564102 168618 588222 169174
rect 588778 168618 588810 169174
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 164898 -2934 165454
rect -2378 164898 19826 165454
rect 20382 164898 55826 165454
rect 56382 164898 91826 165454
rect 92382 164898 127826 165454
rect 128382 164898 163826 165454
rect 164382 164898 199826 165454
rect 200382 164898 235826 165454
rect 236382 164898 271826 165454
rect 272382 164898 307826 165454
rect 308382 164898 343826 165454
rect 344382 164898 379826 165454
rect 380382 164898 415826 165454
rect 416382 164898 451826 165454
rect 452382 164898 487826 165454
rect 488382 164898 523826 165454
rect 524382 164898 559826 165454
rect 560382 164898 586302 165454
rect 586858 164898 586890 165454
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158058 -7734 158614
rect -7178 158058 12986 158614
rect 13542 158058 48986 158614
rect 49542 158058 84986 158614
rect 85542 158058 120986 158614
rect 121542 158058 156986 158614
rect 157542 158058 192986 158614
rect 193542 158058 228986 158614
rect 229542 158058 264986 158614
rect 265542 158058 300986 158614
rect 301542 158058 336986 158614
rect 337542 158058 372986 158614
rect 373542 158058 408986 158614
rect 409542 158058 444986 158614
rect 445542 158058 480986 158614
rect 481542 158058 516986 158614
rect 517542 158058 552986 158614
rect 553542 158058 591102 158614
rect 591658 158058 592650 158614
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154338 -5814 154894
rect -5258 154338 9266 154894
rect 9822 154338 45266 154894
rect 45822 154338 81266 154894
rect 81822 154338 117266 154894
rect 117822 154338 153266 154894
rect 153822 154338 189266 154894
rect 189822 154338 225266 154894
rect 225822 154338 261266 154894
rect 261822 154338 297266 154894
rect 297822 154338 333266 154894
rect 333822 154338 369266 154894
rect 369822 154338 405266 154894
rect 405822 154338 441266 154894
rect 441822 154338 477266 154894
rect 477822 154338 513266 154894
rect 513822 154338 549266 154894
rect 549822 154338 589182 154894
rect 589738 154338 590730 154894
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150618 -3894 151174
rect -3338 150618 5546 151174
rect 6102 150618 41546 151174
rect 42102 150618 77546 151174
rect 78102 150618 113546 151174
rect 114102 150618 149546 151174
rect 150102 150618 185546 151174
rect 186102 150618 221546 151174
rect 222102 150618 257546 151174
rect 258102 150618 293546 151174
rect 294102 150618 329546 151174
rect 330102 150618 365546 151174
rect 366102 150618 401546 151174
rect 402102 150618 437546 151174
rect 438102 150618 473546 151174
rect 474102 150618 509546 151174
rect 510102 150618 545546 151174
rect 546102 150618 581546 151174
rect 582102 150618 587262 151174
rect 587818 150618 588810 151174
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 146898 -1974 147454
rect -1418 146898 1826 147454
rect 2382 146898 37826 147454
rect 38382 146898 73826 147454
rect 74382 146898 109826 147454
rect 110382 146898 145826 147454
rect 146382 146898 181826 147454
rect 182382 146898 217826 147454
rect 218382 146898 253826 147454
rect 254382 146898 289826 147454
rect 290382 146898 325826 147454
rect 326382 146898 361826 147454
rect 362382 146898 397826 147454
rect 398382 146898 433826 147454
rect 434382 146898 469826 147454
rect 470382 146898 505826 147454
rect 506382 146898 541826 147454
rect 542382 146898 577826 147454
rect 578382 146898 585342 147454
rect 585898 146898 586890 147454
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140058 -8694 140614
rect -8138 140058 30986 140614
rect 31542 140058 66986 140614
rect 67542 140058 102986 140614
rect 103542 140058 138986 140614
rect 139542 140058 174986 140614
rect 175542 140058 210986 140614
rect 211542 140058 246986 140614
rect 247542 140058 282986 140614
rect 283542 140058 318986 140614
rect 319542 140058 354986 140614
rect 355542 140058 390986 140614
rect 391542 140058 426986 140614
rect 427542 140058 462986 140614
rect 463542 140058 498986 140614
rect 499542 140058 534986 140614
rect 535542 140058 570986 140614
rect 571542 140058 592062 140614
rect 592618 140058 592650 140614
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136338 -6774 136894
rect -6218 136338 27266 136894
rect 27822 136338 63266 136894
rect 63822 136338 99266 136894
rect 99822 136338 135266 136894
rect 135822 136338 171266 136894
rect 171822 136338 207266 136894
rect 207822 136338 243266 136894
rect 243822 136338 279266 136894
rect 279822 136338 315266 136894
rect 315822 136338 351266 136894
rect 351822 136338 387266 136894
rect 387822 136338 423266 136894
rect 423822 136338 459266 136894
rect 459822 136338 495266 136894
rect 495822 136338 531266 136894
rect 531822 136338 567266 136894
rect 567822 136338 590142 136894
rect 590698 136338 590730 136894
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132618 -4854 133174
rect -4298 132618 23546 133174
rect 24102 132618 59546 133174
rect 60102 132618 95546 133174
rect 96102 132618 131546 133174
rect 132102 132618 167546 133174
rect 168102 132618 203546 133174
rect 204102 132618 239546 133174
rect 240102 132618 275546 133174
rect 276102 132618 311546 133174
rect 312102 132618 347546 133174
rect 348102 132618 383546 133174
rect 384102 132618 419546 133174
rect 420102 132618 455546 133174
rect 456102 132618 491546 133174
rect 492102 132618 527546 133174
rect 528102 132618 563546 133174
rect 564102 132618 588222 133174
rect 588778 132618 588810 133174
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 128898 -2934 129454
rect -2378 128898 19826 129454
rect 20382 128898 55826 129454
rect 56382 128898 91826 129454
rect 92382 128898 127826 129454
rect 128382 128898 163826 129454
rect 164382 128898 199826 129454
rect 200382 128898 235826 129454
rect 236382 128898 271826 129454
rect 272382 128898 307826 129454
rect 308382 128898 343826 129454
rect 344382 128898 379826 129454
rect 380382 128898 415826 129454
rect 416382 128898 451826 129454
rect 452382 128898 487826 129454
rect 488382 128898 523826 129454
rect 524382 128898 559826 129454
rect 560382 128898 586302 129454
rect 586858 128898 586890 129454
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122058 -7734 122614
rect -7178 122058 12986 122614
rect 13542 122058 48986 122614
rect 49542 122058 84986 122614
rect 85542 122058 120986 122614
rect 121542 122058 156986 122614
rect 157542 122058 192986 122614
rect 193542 122058 228986 122614
rect 229542 122058 264986 122614
rect 265542 122058 300986 122614
rect 301542 122058 336986 122614
rect 337542 122058 372986 122614
rect 373542 122058 408986 122614
rect 409542 122058 444986 122614
rect 445542 122058 480986 122614
rect 481542 122058 516986 122614
rect 517542 122058 552986 122614
rect 553542 122058 591102 122614
rect 591658 122058 592650 122614
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118338 -5814 118894
rect -5258 118338 9266 118894
rect 9822 118338 45266 118894
rect 45822 118338 81266 118894
rect 81822 118338 117266 118894
rect 117822 118338 153266 118894
rect 153822 118338 189266 118894
rect 189822 118338 225266 118894
rect 225822 118338 261266 118894
rect 261822 118338 297266 118894
rect 297822 118338 333266 118894
rect 333822 118338 369266 118894
rect 369822 118338 405266 118894
rect 405822 118338 441266 118894
rect 441822 118338 477266 118894
rect 477822 118338 513266 118894
rect 513822 118338 549266 118894
rect 549822 118338 589182 118894
rect 589738 118338 590730 118894
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114618 -3894 115174
rect -3338 114618 5546 115174
rect 6102 114618 41546 115174
rect 42102 114618 77546 115174
rect 78102 114618 113546 115174
rect 114102 114618 149546 115174
rect 150102 114618 185546 115174
rect 186102 114618 221546 115174
rect 222102 114618 257546 115174
rect 258102 114618 293546 115174
rect 294102 114618 329546 115174
rect 330102 114618 365546 115174
rect 366102 114618 401546 115174
rect 402102 114618 437546 115174
rect 438102 114618 473546 115174
rect 474102 114618 509546 115174
rect 510102 114618 545546 115174
rect 546102 114618 581546 115174
rect 582102 114618 587262 115174
rect 587818 114618 588810 115174
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 110898 -1974 111454
rect -1418 110898 1826 111454
rect 2382 110898 37826 111454
rect 38382 110898 73826 111454
rect 74382 110898 109826 111454
rect 110382 110898 145826 111454
rect 146382 110898 181826 111454
rect 182382 110898 217826 111454
rect 218382 110898 253826 111454
rect 254382 110898 289826 111454
rect 290382 110898 325826 111454
rect 326382 110898 361826 111454
rect 362382 110898 397826 111454
rect 398382 110898 433826 111454
rect 434382 110898 469826 111454
rect 470382 110898 505826 111454
rect 506382 110898 541826 111454
rect 542382 110898 577826 111454
rect 578382 110898 585342 111454
rect 585898 110898 586890 111454
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104058 -8694 104614
rect -8138 104058 30986 104614
rect 31542 104058 66986 104614
rect 67542 104058 102986 104614
rect 103542 104058 138986 104614
rect 139542 104058 174986 104614
rect 175542 104058 210986 104614
rect 211542 104058 246986 104614
rect 247542 104058 282986 104614
rect 283542 104058 318986 104614
rect 319542 104058 354986 104614
rect 355542 104058 390986 104614
rect 391542 104058 426986 104614
rect 427542 104058 462986 104614
rect 463542 104058 498986 104614
rect 499542 104058 534986 104614
rect 535542 104058 570986 104614
rect 571542 104058 592062 104614
rect 592618 104058 592650 104614
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100338 -6774 100894
rect -6218 100338 27266 100894
rect 27822 100338 63266 100894
rect 63822 100338 99266 100894
rect 99822 100338 135266 100894
rect 135822 100338 171266 100894
rect 171822 100338 207266 100894
rect 207822 100338 243266 100894
rect 243822 100338 279266 100894
rect 279822 100338 315266 100894
rect 315822 100338 351266 100894
rect 351822 100338 387266 100894
rect 387822 100338 423266 100894
rect 423822 100338 459266 100894
rect 459822 100338 495266 100894
rect 495822 100338 531266 100894
rect 531822 100338 567266 100894
rect 567822 100338 590142 100894
rect 590698 100338 590730 100894
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96618 -4854 97174
rect -4298 96618 23546 97174
rect 24102 96618 59546 97174
rect 60102 96618 95546 97174
rect 96102 96618 131546 97174
rect 132102 96618 167546 97174
rect 168102 96618 203546 97174
rect 204102 96618 239546 97174
rect 240102 96618 275546 97174
rect 276102 96618 311546 97174
rect 312102 96618 347546 97174
rect 348102 96618 383546 97174
rect 384102 96618 419546 97174
rect 420102 96618 455546 97174
rect 456102 96618 491546 97174
rect 492102 96618 527546 97174
rect 528102 96618 563546 97174
rect 564102 96618 588222 97174
rect 588778 96618 588810 97174
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 92898 -2934 93454
rect -2378 92898 19826 93454
rect 20382 92898 55826 93454
rect 56382 92898 91826 93454
rect 92382 92898 127826 93454
rect 128382 92898 163826 93454
rect 164382 92898 199826 93454
rect 200382 92898 235826 93454
rect 236382 92898 271826 93454
rect 272382 92898 307826 93454
rect 308382 92898 343826 93454
rect 344382 92898 379826 93454
rect 380382 92898 415826 93454
rect 416382 92898 451826 93454
rect 452382 92898 487826 93454
rect 488382 92898 523826 93454
rect 524382 92898 559826 93454
rect 560382 92898 586302 93454
rect 586858 92898 586890 93454
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86058 -7734 86614
rect -7178 86058 12986 86614
rect 13542 86058 48986 86614
rect 49542 86058 84986 86614
rect 85542 86058 120986 86614
rect 121542 86058 156986 86614
rect 157542 86058 192986 86614
rect 193542 86058 228986 86614
rect 229542 86058 264986 86614
rect 265542 86058 300986 86614
rect 301542 86058 336986 86614
rect 337542 86058 372986 86614
rect 373542 86058 408986 86614
rect 409542 86058 444986 86614
rect 445542 86058 480986 86614
rect 481542 86058 516986 86614
rect 517542 86058 552986 86614
rect 553542 86058 591102 86614
rect 591658 86058 592650 86614
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82338 -5814 82894
rect -5258 82338 9266 82894
rect 9822 82338 45266 82894
rect 45822 82338 81266 82894
rect 81822 82338 117266 82894
rect 117822 82338 153266 82894
rect 153822 82338 189266 82894
rect 189822 82338 225266 82894
rect 225822 82338 261266 82894
rect 261822 82338 297266 82894
rect 297822 82338 333266 82894
rect 333822 82338 369266 82894
rect 369822 82338 405266 82894
rect 405822 82338 441266 82894
rect 441822 82338 477266 82894
rect 477822 82338 513266 82894
rect 513822 82338 549266 82894
rect 549822 82338 589182 82894
rect 589738 82338 590730 82894
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78618 -3894 79174
rect -3338 78618 5546 79174
rect 6102 78618 41546 79174
rect 42102 78618 77546 79174
rect 78102 78618 113546 79174
rect 114102 78618 149546 79174
rect 150102 78618 185546 79174
rect 186102 78618 221546 79174
rect 222102 78618 257546 79174
rect 258102 78618 293546 79174
rect 294102 78618 329546 79174
rect 330102 78618 365546 79174
rect 366102 78618 401546 79174
rect 402102 78618 437546 79174
rect 438102 78618 473546 79174
rect 474102 78618 509546 79174
rect 510102 78618 545546 79174
rect 546102 78618 581546 79174
rect 582102 78618 587262 79174
rect 587818 78618 588810 79174
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 74898 -1974 75454
rect -1418 74898 1826 75454
rect 2382 74898 37826 75454
rect 38382 74898 73826 75454
rect 74382 74898 109826 75454
rect 110382 74898 145826 75454
rect 146382 74898 181826 75454
rect 182382 74898 217826 75454
rect 218382 74898 253826 75454
rect 254382 74898 289826 75454
rect 290382 74898 325826 75454
rect 326382 74898 361826 75454
rect 362382 74898 397826 75454
rect 398382 74898 433826 75454
rect 434382 74898 469826 75454
rect 470382 74898 505826 75454
rect 506382 74898 541826 75454
rect 542382 74898 577826 75454
rect 578382 74898 585342 75454
rect 585898 74898 586890 75454
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68058 -8694 68614
rect -8138 68058 30986 68614
rect 31542 68058 66986 68614
rect 67542 68058 102986 68614
rect 103542 68058 138986 68614
rect 139542 68058 174986 68614
rect 175542 68058 210986 68614
rect 211542 68058 246986 68614
rect 247542 68058 282986 68614
rect 283542 68058 318986 68614
rect 319542 68058 354986 68614
rect 355542 68058 390986 68614
rect 391542 68058 426986 68614
rect 427542 68058 462986 68614
rect 463542 68058 498986 68614
rect 499542 68058 534986 68614
rect 535542 68058 570986 68614
rect 571542 68058 592062 68614
rect 592618 68058 592650 68614
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64338 -6774 64894
rect -6218 64338 27266 64894
rect 27822 64338 63266 64894
rect 63822 64338 99266 64894
rect 99822 64338 135266 64894
rect 135822 64338 171266 64894
rect 171822 64338 207266 64894
rect 207822 64338 243266 64894
rect 243822 64338 279266 64894
rect 279822 64338 315266 64894
rect 315822 64338 351266 64894
rect 351822 64338 387266 64894
rect 387822 64338 423266 64894
rect 423822 64338 459266 64894
rect 459822 64338 495266 64894
rect 495822 64338 531266 64894
rect 531822 64338 567266 64894
rect 567822 64338 590142 64894
rect 590698 64338 590730 64894
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60618 -4854 61174
rect -4298 60618 23546 61174
rect 24102 60618 59546 61174
rect 60102 60618 95546 61174
rect 96102 60618 131546 61174
rect 132102 60618 167546 61174
rect 168102 60618 203546 61174
rect 204102 60618 239546 61174
rect 240102 60618 275546 61174
rect 276102 60618 311546 61174
rect 312102 60618 347546 61174
rect 348102 60618 383546 61174
rect 384102 60618 419546 61174
rect 420102 60618 455546 61174
rect 456102 60618 491546 61174
rect 492102 60618 527546 61174
rect 528102 60618 563546 61174
rect 564102 60618 588222 61174
rect 588778 60618 588810 61174
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 56898 -2934 57454
rect -2378 56898 19826 57454
rect 20382 56898 55826 57454
rect 56382 56898 91826 57454
rect 92382 56898 127826 57454
rect 128382 56898 163826 57454
rect 164382 56898 199826 57454
rect 200382 56898 235826 57454
rect 236382 56898 271826 57454
rect 272382 56898 307826 57454
rect 308382 56898 343826 57454
rect 344382 56898 379826 57454
rect 380382 56898 415826 57454
rect 416382 56898 451826 57454
rect 452382 56898 487826 57454
rect 488382 56898 523826 57454
rect 524382 56898 559826 57454
rect 560382 56898 586302 57454
rect 586858 56898 586890 57454
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50058 -7734 50614
rect -7178 50058 12986 50614
rect 13542 50058 48986 50614
rect 49542 50058 84986 50614
rect 85542 50058 120986 50614
rect 121542 50058 156986 50614
rect 157542 50058 192986 50614
rect 193542 50058 228986 50614
rect 229542 50058 264986 50614
rect 265542 50058 300986 50614
rect 301542 50058 336986 50614
rect 337542 50058 372986 50614
rect 373542 50058 408986 50614
rect 409542 50058 444986 50614
rect 445542 50058 480986 50614
rect 481542 50058 516986 50614
rect 517542 50058 552986 50614
rect 553542 50058 591102 50614
rect 591658 50058 592650 50614
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46338 -5814 46894
rect -5258 46338 9266 46894
rect 9822 46338 45266 46894
rect 45822 46338 81266 46894
rect 81822 46338 117266 46894
rect 117822 46338 153266 46894
rect 153822 46338 189266 46894
rect 189822 46338 225266 46894
rect 225822 46338 261266 46894
rect 261822 46338 297266 46894
rect 297822 46338 333266 46894
rect 333822 46338 369266 46894
rect 369822 46338 405266 46894
rect 405822 46338 441266 46894
rect 441822 46338 477266 46894
rect 477822 46338 513266 46894
rect 513822 46338 549266 46894
rect 549822 46338 589182 46894
rect 589738 46338 590730 46894
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42618 -3894 43174
rect -3338 42618 5546 43174
rect 6102 42618 41546 43174
rect 42102 42618 77546 43174
rect 78102 42618 113546 43174
rect 114102 42618 149546 43174
rect 150102 42618 185546 43174
rect 186102 42618 221546 43174
rect 222102 42618 257546 43174
rect 258102 42618 293546 43174
rect 294102 42618 329546 43174
rect 330102 42618 365546 43174
rect 366102 42618 401546 43174
rect 402102 42618 437546 43174
rect 438102 42618 473546 43174
rect 474102 42618 509546 43174
rect 510102 42618 545546 43174
rect 546102 42618 581546 43174
rect 582102 42618 587262 43174
rect 587818 42618 588810 43174
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 38898 -1974 39454
rect -1418 38898 1826 39454
rect 2382 38898 37826 39454
rect 38382 38898 73826 39454
rect 74382 38898 109826 39454
rect 110382 38898 145826 39454
rect 146382 38898 181826 39454
rect 182382 38898 217826 39454
rect 218382 38898 253826 39454
rect 254382 38898 289826 39454
rect 290382 38898 325826 39454
rect 326382 38898 361826 39454
rect 362382 38898 397826 39454
rect 398382 38898 433826 39454
rect 434382 38898 469826 39454
rect 470382 38898 505826 39454
rect 506382 38898 541826 39454
rect 542382 38898 577826 39454
rect 578382 38898 585342 39454
rect 585898 38898 586890 39454
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32058 -8694 32614
rect -8138 32058 30986 32614
rect 31542 32058 66986 32614
rect 67542 32058 102986 32614
rect 103542 32058 138986 32614
rect 139542 32058 174986 32614
rect 175542 32058 210986 32614
rect 211542 32058 246986 32614
rect 247542 32058 282986 32614
rect 283542 32058 318986 32614
rect 319542 32058 354986 32614
rect 355542 32058 390986 32614
rect 391542 32058 426986 32614
rect 427542 32058 462986 32614
rect 463542 32058 498986 32614
rect 499542 32058 534986 32614
rect 535542 32058 570986 32614
rect 571542 32058 592062 32614
rect 592618 32058 592650 32614
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28338 -6774 28894
rect -6218 28338 27266 28894
rect 27822 28338 63266 28894
rect 63822 28338 99266 28894
rect 99822 28338 135266 28894
rect 135822 28338 171266 28894
rect 171822 28338 207266 28894
rect 207822 28338 243266 28894
rect 243822 28338 279266 28894
rect 279822 28338 315266 28894
rect 315822 28338 351266 28894
rect 351822 28338 387266 28894
rect 387822 28338 423266 28894
rect 423822 28338 459266 28894
rect 459822 28338 495266 28894
rect 495822 28338 531266 28894
rect 531822 28338 567266 28894
rect 567822 28338 590142 28894
rect 590698 28338 590730 28894
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24618 -4854 25174
rect -4298 24618 23546 25174
rect 24102 24618 59546 25174
rect 60102 24618 95546 25174
rect 96102 24618 131546 25174
rect 132102 24618 167546 25174
rect 168102 24618 203546 25174
rect 204102 24618 239546 25174
rect 240102 24618 275546 25174
rect 276102 24618 311546 25174
rect 312102 24618 347546 25174
rect 348102 24618 383546 25174
rect 384102 24618 419546 25174
rect 420102 24618 455546 25174
rect 456102 24618 491546 25174
rect 492102 24618 527546 25174
rect 528102 24618 563546 25174
rect 564102 24618 588222 25174
rect 588778 24618 588810 25174
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 20898 -2934 21454
rect -2378 20898 19826 21454
rect 20382 20898 55826 21454
rect 56382 20898 91826 21454
rect 92382 20898 127826 21454
rect 128382 20898 163826 21454
rect 164382 20898 199826 21454
rect 200382 20898 235826 21454
rect 236382 20898 271826 21454
rect 272382 20898 307826 21454
rect 308382 20898 343826 21454
rect 344382 20898 379826 21454
rect 380382 20898 415826 21454
rect 416382 20898 451826 21454
rect 452382 20898 487826 21454
rect 488382 20898 523826 21454
rect 524382 20898 559826 21454
rect 560382 20898 586302 21454
rect 586858 20898 586890 21454
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14058 -7734 14614
rect -7178 14058 12986 14614
rect 13542 14058 48986 14614
rect 49542 14058 84986 14614
rect 85542 14058 120986 14614
rect 121542 14058 156986 14614
rect 157542 14058 192986 14614
rect 193542 14058 228986 14614
rect 229542 14058 264986 14614
rect 265542 14058 300986 14614
rect 301542 14058 336986 14614
rect 337542 14058 372986 14614
rect 373542 14058 408986 14614
rect 409542 14058 444986 14614
rect 445542 14058 480986 14614
rect 481542 14058 516986 14614
rect 517542 14058 552986 14614
rect 553542 14058 591102 14614
rect 591658 14058 592650 14614
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10338 -5814 10894
rect -5258 10338 9266 10894
rect 9822 10338 45266 10894
rect 45822 10338 81266 10894
rect 81822 10338 117266 10894
rect 117822 10338 153266 10894
rect 153822 10338 189266 10894
rect 189822 10338 225266 10894
rect 225822 10338 261266 10894
rect 261822 10338 297266 10894
rect 297822 10338 333266 10894
rect 333822 10338 369266 10894
rect 369822 10338 405266 10894
rect 405822 10338 441266 10894
rect 441822 10338 477266 10894
rect 477822 10338 513266 10894
rect 513822 10338 549266 10894
rect 549822 10338 589182 10894
rect 589738 10338 590730 10894
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6618 -3894 7174
rect -3338 6618 5546 7174
rect 6102 6618 41546 7174
rect 42102 6618 77546 7174
rect 78102 6618 113546 7174
rect 114102 6618 149546 7174
rect 150102 6618 185546 7174
rect 186102 6618 221546 7174
rect 222102 6618 257546 7174
rect 258102 6618 293546 7174
rect 294102 6618 329546 7174
rect 330102 6618 365546 7174
rect 366102 6618 401546 7174
rect 402102 6618 437546 7174
rect 438102 6618 473546 7174
rect 474102 6618 509546 7174
rect 510102 6618 545546 7174
rect 546102 6618 581546 7174
rect 582102 6618 587262 7174
rect 587818 6618 588810 7174
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 2898 -1974 3454
rect -1418 2898 1826 3454
rect 2382 2898 37826 3454
rect 38382 2898 73826 3454
rect 74382 2898 109826 3454
rect 110382 2898 145826 3454
rect 146382 2898 181826 3454
rect 182382 2898 217826 3454
rect 218382 2898 253826 3454
rect 254382 2898 289826 3454
rect 290382 2898 325826 3454
rect 326382 2898 361826 3454
rect 362382 2898 397826 3454
rect 398382 2898 433826 3454
rect 434382 2898 469826 3454
rect 470382 2898 505826 3454
rect 506382 2898 541826 3454
rect 542382 2898 577826 3454
rect 578382 2898 585342 3454
rect 585898 2898 586890 3454
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -902 -1974 -346
rect -1418 -902 1826 -346
rect 2382 -902 37826 -346
rect 38382 -902 73826 -346
rect 74382 -902 109826 -346
rect 110382 -902 145826 -346
rect 146382 -902 181826 -346
rect 182382 -902 217826 -346
rect 218382 -902 253826 -346
rect 254382 -902 289826 -346
rect 290382 -902 325826 -346
rect 326382 -902 361826 -346
rect 362382 -902 397826 -346
rect 398382 -902 433826 -346
rect 434382 -902 469826 -346
rect 470382 -902 505826 -346
rect 506382 -902 541826 -346
rect 542382 -902 577826 -346
rect 578382 -902 585342 -346
rect 585898 -902 585930 -346
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1862 -2934 -1306
rect -2378 -1862 19826 -1306
rect 20382 -1862 55826 -1306
rect 56382 -1862 91826 -1306
rect 92382 -1862 127826 -1306
rect 128382 -1862 163826 -1306
rect 164382 -1862 199826 -1306
rect 200382 -1862 235826 -1306
rect 236382 -1862 271826 -1306
rect 272382 -1862 307826 -1306
rect 308382 -1862 343826 -1306
rect 344382 -1862 379826 -1306
rect 380382 -1862 415826 -1306
rect 416382 -1862 451826 -1306
rect 452382 -1862 487826 -1306
rect 488382 -1862 523826 -1306
rect 524382 -1862 559826 -1306
rect 560382 -1862 586302 -1306
rect 586858 -1862 586890 -1306
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2822 -3894 -2266
rect -3338 -2822 5546 -2266
rect 6102 -2822 41546 -2266
rect 42102 -2822 77546 -2266
rect 78102 -2822 113546 -2266
rect 114102 -2822 149546 -2266
rect 150102 -2822 185546 -2266
rect 186102 -2822 221546 -2266
rect 222102 -2822 257546 -2266
rect 258102 -2822 293546 -2266
rect 294102 -2822 329546 -2266
rect 330102 -2822 365546 -2266
rect 366102 -2822 401546 -2266
rect 402102 -2822 437546 -2266
rect 438102 -2822 473546 -2266
rect 474102 -2822 509546 -2266
rect 510102 -2822 545546 -2266
rect 546102 -2822 581546 -2266
rect 582102 -2822 587262 -2266
rect 587818 -2822 587850 -2266
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3782 -4854 -3226
rect -4298 -3782 23546 -3226
rect 24102 -3782 59546 -3226
rect 60102 -3782 95546 -3226
rect 96102 -3782 131546 -3226
rect 132102 -3782 167546 -3226
rect 168102 -3782 203546 -3226
rect 204102 -3782 239546 -3226
rect 240102 -3782 275546 -3226
rect 276102 -3782 311546 -3226
rect 312102 -3782 347546 -3226
rect 348102 -3782 383546 -3226
rect 384102 -3782 419546 -3226
rect 420102 -3782 455546 -3226
rect 456102 -3782 491546 -3226
rect 492102 -3782 527546 -3226
rect 528102 -3782 563546 -3226
rect 564102 -3782 588222 -3226
rect 588778 -3782 588810 -3226
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4742 -5814 -4186
rect -5258 -4742 9266 -4186
rect 9822 -4742 45266 -4186
rect 45822 -4742 81266 -4186
rect 81822 -4742 117266 -4186
rect 117822 -4742 153266 -4186
rect 153822 -4742 189266 -4186
rect 189822 -4742 225266 -4186
rect 225822 -4742 261266 -4186
rect 261822 -4742 297266 -4186
rect 297822 -4742 333266 -4186
rect 333822 -4742 369266 -4186
rect 369822 -4742 405266 -4186
rect 405822 -4742 441266 -4186
rect 441822 -4742 477266 -4186
rect 477822 -4742 513266 -4186
rect 513822 -4742 549266 -4186
rect 549822 -4742 589182 -4186
rect 589738 -4742 589770 -4186
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5702 -6774 -5146
rect -6218 -5702 27266 -5146
rect 27822 -5702 63266 -5146
rect 63822 -5702 99266 -5146
rect 99822 -5702 135266 -5146
rect 135822 -5702 171266 -5146
rect 171822 -5702 207266 -5146
rect 207822 -5702 243266 -5146
rect 243822 -5702 279266 -5146
rect 279822 -5702 315266 -5146
rect 315822 -5702 351266 -5146
rect 351822 -5702 387266 -5146
rect 387822 -5702 423266 -5146
rect 423822 -5702 459266 -5146
rect 459822 -5702 495266 -5146
rect 495822 -5702 531266 -5146
rect 531822 -5702 567266 -5146
rect 567822 -5702 590142 -5146
rect 590698 -5702 590730 -5146
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6662 -7734 -6106
rect -7178 -6662 12986 -6106
rect 13542 -6662 48986 -6106
rect 49542 -6662 84986 -6106
rect 85542 -6662 120986 -6106
rect 121542 -6662 156986 -6106
rect 157542 -6662 192986 -6106
rect 193542 -6662 228986 -6106
rect 229542 -6662 264986 -6106
rect 265542 -6662 300986 -6106
rect 301542 -6662 336986 -6106
rect 337542 -6662 372986 -6106
rect 373542 -6662 408986 -6106
rect 409542 -6662 444986 -6106
rect 445542 -6662 480986 -6106
rect 481542 -6662 516986 -6106
rect 517542 -6662 552986 -6106
rect 553542 -6662 591102 -6106
rect 591658 -6662 591690 -6106
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7622 -8694 -7066
rect -8138 -7622 30986 -7066
rect 31542 -7622 66986 -7066
rect 67542 -7622 102986 -7066
rect 103542 -7622 138986 -7066
rect 139542 -7622 174986 -7066
rect 175542 -7622 210986 -7066
rect 211542 -7622 246986 -7066
rect 247542 -7622 282986 -7066
rect 283542 -7622 318986 -7066
rect 319542 -7622 354986 -7066
rect 355542 -7622 390986 -7066
rect 391542 -7622 426986 -7066
rect 427542 -7622 462986 -7066
rect 463542 -7622 498986 -7066
rect 499542 -7622 534986 -7066
rect 535542 -7622 570986 -7066
rect 571542 -7622 592062 -7066
rect 592618 -7622 592650 -7066
rect -8726 -7654 592650 -7622
use user_proj_example  mprj
timestamp 1634570663
transform 1 0 235000 0 1 338000
box 18 0 59878 40000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 4 analog_io[0]
port 1 nsew
rlabel metal2 s 446098 703520 446210 704960 4 analog_io[10]
port 2 nsew
rlabel metal2 s 381146 703520 381258 704960 4 analog_io[11]
port 3 nsew
rlabel metal2 s 316286 703520 316398 704960 4 analog_io[12]
port 4 nsew
rlabel metal2 s 251426 703520 251538 704960 4 analog_io[13]
port 5 nsew
rlabel metal2 s 186474 703520 186586 704960 4 analog_io[14]
port 6 nsew
rlabel metal2 s 121614 703520 121726 704960 4 analog_io[15]
port 7 nsew
rlabel metal2 s 56754 703520 56866 704960 4 analog_io[16]
port 8 nsew
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 9 nsew
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 10 nsew
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 11 nsew
rlabel metal3 s 583520 338452 584960 338692 4 analog_io[1]
port 12 nsew
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 13 nsew
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 14 nsew
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 15 nsew
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 16 nsew
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 17 nsew
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 18 nsew
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 19 nsew
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 20 nsew
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 21 nsew
rlabel metal3 s 583520 391628 584960 391868 4 analog_io[2]
port 22 nsew
rlabel metal3 s 583520 444668 584960 444908 4 analog_io[3]
port 23 nsew
rlabel metal3 s 583520 497844 584960 498084 4 analog_io[4]
port 24 nsew
rlabel metal3 s 583520 551020 584960 551260 4 analog_io[5]
port 25 nsew
rlabel metal3 s 583520 604060 584960 604300 4 analog_io[6]
port 26 nsew
rlabel metal3 s 583520 657236 584960 657476 4 analog_io[7]
port 27 nsew
rlabel metal2 s 575818 703520 575930 704960 4 analog_io[8]
port 28 nsew
rlabel metal2 s 510958 703520 511070 704960 4 analog_io[9]
port 29 nsew
rlabel metal3 s 583520 6476 584960 6716 4 io_in[0]
port 30 nsew
rlabel metal3 s 583520 457996 584960 458236 4 io_in[10]
port 31 nsew
rlabel metal3 s 583520 511172 584960 511412 4 io_in[11]
port 32 nsew
rlabel metal3 s 583520 564212 584960 564452 4 io_in[12]
port 33 nsew
rlabel metal3 s 583520 617388 584960 617628 4 io_in[13]
port 34 nsew
rlabel metal3 s 583520 670564 584960 670804 4 io_in[14]
port 35 nsew
rlabel metal2 s 559626 703520 559738 704960 4 io_in[15]
port 36 nsew
rlabel metal2 s 494766 703520 494878 704960 4 io_in[16]
port 37 nsew
rlabel metal2 s 429814 703520 429926 704960 4 io_in[17]
port 38 nsew
rlabel metal2 s 364954 703520 365066 704960 4 io_in[18]
port 39 nsew
rlabel metal2 s 300094 703520 300206 704960 4 io_in[19]
port 40 nsew
rlabel metal3 s 583520 46188 584960 46428 4 io_in[1]
port 41 nsew
rlabel metal2 s 235142 703520 235254 704960 4 io_in[20]
port 42 nsew
rlabel metal2 s 170282 703520 170394 704960 4 io_in[21]
port 43 nsew
rlabel metal2 s 105422 703520 105534 704960 4 io_in[22]
port 44 nsew
rlabel metal2 s 40470 703520 40582 704960 4 io_in[23]
port 45 nsew
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 46 nsew
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 47 nsew
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 48 nsew
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 49 nsew
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 50 nsew
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 51 nsew
rlabel metal3 s 583520 86036 584960 86276 4 io_in[2]
port 52 nsew
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 53 nsew
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 54 nsew
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 55 nsew
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 56 nsew
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 57 nsew
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 58 nsew
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 59 nsew
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 60 nsew
rlabel metal3 s 583520 125884 584960 126124 4 io_in[3]
port 61 nsew
rlabel metal3 s 583520 165732 584960 165972 4 io_in[4]
port 62 nsew
rlabel metal3 s 583520 205580 584960 205820 4 io_in[5]
port 63 nsew
rlabel metal3 s 583520 245428 584960 245668 4 io_in[6]
port 64 nsew
rlabel metal3 s 583520 298604 584960 298844 4 io_in[7]
port 65 nsew
rlabel metal3 s 583520 351780 584960 352020 4 io_in[8]
port 66 nsew
rlabel metal3 s 583520 404820 584960 405060 4 io_in[9]
port 67 nsew
rlabel metal3 s 583520 32996 584960 33236 4 io_oeb[0]
port 68 nsew
rlabel metal3 s 583520 484516 584960 484756 4 io_oeb[10]
port 69 nsew
rlabel metal3 s 583520 537692 584960 537932 4 io_oeb[11]
port 70 nsew
rlabel metal3 s 583520 590868 584960 591108 4 io_oeb[12]
port 71 nsew
rlabel metal3 s 583520 643908 584960 644148 4 io_oeb[13]
port 72 nsew
rlabel metal3 s 583520 697084 584960 697324 4 io_oeb[14]
port 73 nsew
rlabel metal2 s 527150 703520 527262 704960 4 io_oeb[15]
port 74 nsew
rlabel metal2 s 462290 703520 462402 704960 4 io_oeb[16]
port 75 nsew
rlabel metal2 s 397430 703520 397542 704960 4 io_oeb[17]
port 76 nsew
rlabel metal2 s 332478 703520 332590 704960 4 io_oeb[18]
port 77 nsew
rlabel metal2 s 267618 703520 267730 704960 4 io_oeb[19]
port 78 nsew
rlabel metal3 s 583520 72844 584960 73084 4 io_oeb[1]
port 79 nsew
rlabel metal2 s 202758 703520 202870 704960 4 io_oeb[20]
port 80 nsew
rlabel metal2 s 137806 703520 137918 704960 4 io_oeb[21]
port 81 nsew
rlabel metal2 s 72946 703520 73058 704960 4 io_oeb[22]
port 82 nsew
rlabel metal2 s 8086 703520 8198 704960 4 io_oeb[23]
port 83 nsew
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 84 nsew
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 85 nsew
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 86 nsew
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 87 nsew
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 88 nsew
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 89 nsew
rlabel metal3 s 583520 112692 584960 112932 4 io_oeb[2]
port 90 nsew
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 91 nsew
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 92 nsew
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 93 nsew
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 94 nsew
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 95 nsew
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 96 nsew
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 97 nsew
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 98 nsew
rlabel metal3 s 583520 152540 584960 152780 4 io_oeb[3]
port 99 nsew
rlabel metal3 s 583520 192388 584960 192628 4 io_oeb[4]
port 100 nsew
rlabel metal3 s 583520 232236 584960 232476 4 io_oeb[5]
port 101 nsew
rlabel metal3 s 583520 272084 584960 272324 4 io_oeb[6]
port 102 nsew
rlabel metal3 s 583520 325124 584960 325364 4 io_oeb[7]
port 103 nsew
rlabel metal3 s 583520 378300 584960 378540 4 io_oeb[8]
port 104 nsew
rlabel metal3 s 583520 431476 584960 431716 4 io_oeb[9]
port 105 nsew
rlabel metal3 s 583520 19668 584960 19908 4 io_out[0]
port 106 nsew
rlabel metal3 s 583520 471324 584960 471564 4 io_out[10]
port 107 nsew
rlabel metal3 s 583520 524364 584960 524604 4 io_out[11]
port 108 nsew
rlabel metal3 s 583520 577540 584960 577780 4 io_out[12]
port 109 nsew
rlabel metal3 s 583520 630716 584960 630956 4 io_out[13]
port 110 nsew
rlabel metal3 s 583520 683756 584960 683996 4 io_out[14]
port 111 nsew
rlabel metal2 s 543434 703520 543546 704960 4 io_out[15]
port 112 nsew
rlabel metal2 s 478482 703520 478594 704960 4 io_out[16]
port 113 nsew
rlabel metal2 s 413622 703520 413734 704960 4 io_out[17]
port 114 nsew
rlabel metal2 s 348762 703520 348874 704960 4 io_out[18]
port 115 nsew
rlabel metal2 s 283810 703520 283922 704960 4 io_out[19]
port 116 nsew
rlabel metal3 s 583520 59516 584960 59756 4 io_out[1]
port 117 nsew
rlabel metal2 s 218950 703520 219062 704960 4 io_out[20]
port 118 nsew
rlabel metal2 s 154090 703520 154202 704960 4 io_out[21]
port 119 nsew
rlabel metal2 s 89138 703520 89250 704960 4 io_out[22]
port 120 nsew
rlabel metal2 s 24278 703520 24390 704960 4 io_out[23]
port 121 nsew
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 122 nsew
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 123 nsew
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 124 nsew
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 125 nsew
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 126 nsew
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 127 nsew
rlabel metal3 s 583520 99364 584960 99604 4 io_out[2]
port 128 nsew
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 129 nsew
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 130 nsew
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 131 nsew
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 132 nsew
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 133 nsew
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 134 nsew
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 135 nsew
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 136 nsew
rlabel metal3 s 583520 139212 584960 139452 4 io_out[3]
port 137 nsew
rlabel metal3 s 583520 179060 584960 179300 4 io_out[4]
port 138 nsew
rlabel metal3 s 583520 218908 584960 219148 4 io_out[5]
port 139 nsew
rlabel metal3 s 583520 258756 584960 258996 4 io_out[6]
port 140 nsew
rlabel metal3 s 583520 311932 584960 312172 4 io_out[7]
port 141 nsew
rlabel metal3 s 583520 364972 584960 365212 4 io_out[8]
port 142 nsew
rlabel metal3 s 583520 418148 584960 418388 4 io_out[9]
port 143 nsew
rlabel metal2 s 125846 -960 125958 480 4 la_data_in[0]
port 144 nsew
rlabel metal2 s 480506 -960 480618 480 4 la_data_in[100]
port 145 nsew
rlabel metal2 s 484002 -960 484114 480 4 la_data_in[101]
port 146 nsew
rlabel metal2 s 487590 -960 487702 480 4 la_data_in[102]
port 147 nsew
rlabel metal2 s 491086 -960 491198 480 4 la_data_in[103]
port 148 nsew
rlabel metal2 s 494674 -960 494786 480 4 la_data_in[104]
port 149 nsew
rlabel metal2 s 498170 -960 498282 480 4 la_data_in[105]
port 150 nsew
rlabel metal2 s 501758 -960 501870 480 4 la_data_in[106]
port 151 nsew
rlabel metal2 s 505346 -960 505458 480 4 la_data_in[107]
port 152 nsew
rlabel metal2 s 508842 -960 508954 480 4 la_data_in[108]
port 153 nsew
rlabel metal2 s 512430 -960 512542 480 4 la_data_in[109]
port 154 nsew
rlabel metal2 s 161266 -960 161378 480 4 la_data_in[10]
port 155 nsew
rlabel metal2 s 515926 -960 516038 480 4 la_data_in[110]
port 156 nsew
rlabel metal2 s 519514 -960 519626 480 4 la_data_in[111]
port 157 nsew
rlabel metal2 s 523010 -960 523122 480 4 la_data_in[112]
port 158 nsew
rlabel metal2 s 526598 -960 526710 480 4 la_data_in[113]
port 159 nsew
rlabel metal2 s 530094 -960 530206 480 4 la_data_in[114]
port 160 nsew
rlabel metal2 s 533682 -960 533794 480 4 la_data_in[115]
port 161 nsew
rlabel metal2 s 537178 -960 537290 480 4 la_data_in[116]
port 162 nsew
rlabel metal2 s 540766 -960 540878 480 4 la_data_in[117]
port 163 nsew
rlabel metal2 s 544354 -960 544466 480 4 la_data_in[118]
port 164 nsew
rlabel metal2 s 547850 -960 547962 480 4 la_data_in[119]
port 165 nsew
rlabel metal2 s 164854 -960 164966 480 4 la_data_in[11]
port 166 nsew
rlabel metal2 s 551438 -960 551550 480 4 la_data_in[120]
port 167 nsew
rlabel metal2 s 554934 -960 555046 480 4 la_data_in[121]
port 168 nsew
rlabel metal2 s 558522 -960 558634 480 4 la_data_in[122]
port 169 nsew
rlabel metal2 s 562018 -960 562130 480 4 la_data_in[123]
port 170 nsew
rlabel metal2 s 565606 -960 565718 480 4 la_data_in[124]
port 171 nsew
rlabel metal2 s 569102 -960 569214 480 4 la_data_in[125]
port 172 nsew
rlabel metal2 s 572690 -960 572802 480 4 la_data_in[126]
port 173 nsew
rlabel metal2 s 576278 -960 576390 480 4 la_data_in[127]
port 174 nsew
rlabel metal2 s 168350 -960 168462 480 4 la_data_in[12]
port 175 nsew
rlabel metal2 s 171938 -960 172050 480 4 la_data_in[13]
port 176 nsew
rlabel metal2 s 175434 -960 175546 480 4 la_data_in[14]
port 177 nsew
rlabel metal2 s 179022 -960 179134 480 4 la_data_in[15]
port 178 nsew
rlabel metal2 s 182518 -960 182630 480 4 la_data_in[16]
port 179 nsew
rlabel metal2 s 186106 -960 186218 480 4 la_data_in[17]
port 180 nsew
rlabel metal2 s 189694 -960 189806 480 4 la_data_in[18]
port 181 nsew
rlabel metal2 s 193190 -960 193302 480 4 la_data_in[19]
port 182 nsew
rlabel metal2 s 129342 -960 129454 480 4 la_data_in[1]
port 183 nsew
rlabel metal2 s 196778 -960 196890 480 4 la_data_in[20]
port 184 nsew
rlabel metal2 s 200274 -960 200386 480 4 la_data_in[21]
port 185 nsew
rlabel metal2 s 203862 -960 203974 480 4 la_data_in[22]
port 186 nsew
rlabel metal2 s 207358 -960 207470 480 4 la_data_in[23]
port 187 nsew
rlabel metal2 s 210946 -960 211058 480 4 la_data_in[24]
port 188 nsew
rlabel metal2 s 214442 -960 214554 480 4 la_data_in[25]
port 189 nsew
rlabel metal2 s 218030 -960 218142 480 4 la_data_in[26]
port 190 nsew
rlabel metal2 s 221526 -960 221638 480 4 la_data_in[27]
port 191 nsew
rlabel metal2 s 225114 -960 225226 480 4 la_data_in[28]
port 192 nsew
rlabel metal2 s 228702 -960 228814 480 4 la_data_in[29]
port 193 nsew
rlabel metal2 s 132930 -960 133042 480 4 la_data_in[2]
port 194 nsew
rlabel metal2 s 232198 -960 232310 480 4 la_data_in[30]
port 195 nsew
rlabel metal2 s 235786 -960 235898 480 4 la_data_in[31]
port 196 nsew
rlabel metal2 s 239282 -960 239394 480 4 la_data_in[32]
port 197 nsew
rlabel metal2 s 242870 -960 242982 480 4 la_data_in[33]
port 198 nsew
rlabel metal2 s 246366 -960 246478 480 4 la_data_in[34]
port 199 nsew
rlabel metal2 s 249954 -960 250066 480 4 la_data_in[35]
port 200 nsew
rlabel metal2 s 253450 -960 253562 480 4 la_data_in[36]
port 201 nsew
rlabel metal2 s 257038 -960 257150 480 4 la_data_in[37]
port 202 nsew
rlabel metal2 s 260626 -960 260738 480 4 la_data_in[38]
port 203 nsew
rlabel metal2 s 264122 -960 264234 480 4 la_data_in[39]
port 204 nsew
rlabel metal2 s 136426 -960 136538 480 4 la_data_in[3]
port 205 nsew
rlabel metal2 s 267710 -960 267822 480 4 la_data_in[40]
port 206 nsew
rlabel metal2 s 271206 -960 271318 480 4 la_data_in[41]
port 207 nsew
rlabel metal2 s 274794 -960 274906 480 4 la_data_in[42]
port 208 nsew
rlabel metal2 s 278290 -960 278402 480 4 la_data_in[43]
port 209 nsew
rlabel metal2 s 281878 -960 281990 480 4 la_data_in[44]
port 210 nsew
rlabel metal2 s 285374 -960 285486 480 4 la_data_in[45]
port 211 nsew
rlabel metal2 s 288962 -960 289074 480 4 la_data_in[46]
port 212 nsew
rlabel metal2 s 292550 -960 292662 480 4 la_data_in[47]
port 213 nsew
rlabel metal2 s 296046 -960 296158 480 4 la_data_in[48]
port 214 nsew
rlabel metal2 s 299634 -960 299746 480 4 la_data_in[49]
port 215 nsew
rlabel metal2 s 140014 -960 140126 480 4 la_data_in[4]
port 216 nsew
rlabel metal2 s 303130 -960 303242 480 4 la_data_in[50]
port 217 nsew
rlabel metal2 s 306718 -960 306830 480 4 la_data_in[51]
port 218 nsew
rlabel metal2 s 310214 -960 310326 480 4 la_data_in[52]
port 219 nsew
rlabel metal2 s 313802 -960 313914 480 4 la_data_in[53]
port 220 nsew
rlabel metal2 s 317298 -960 317410 480 4 la_data_in[54]
port 221 nsew
rlabel metal2 s 320886 -960 320998 480 4 la_data_in[55]
port 222 nsew
rlabel metal2 s 324382 -960 324494 480 4 la_data_in[56]
port 223 nsew
rlabel metal2 s 327970 -960 328082 480 4 la_data_in[57]
port 224 nsew
rlabel metal2 s 331558 -960 331670 480 4 la_data_in[58]
port 225 nsew
rlabel metal2 s 335054 -960 335166 480 4 la_data_in[59]
port 226 nsew
rlabel metal2 s 143510 -960 143622 480 4 la_data_in[5]
port 227 nsew
rlabel metal2 s 338642 -960 338754 480 4 la_data_in[60]
port 228 nsew
rlabel metal2 s 342138 -960 342250 480 4 la_data_in[61]
port 229 nsew
rlabel metal2 s 345726 -960 345838 480 4 la_data_in[62]
port 230 nsew
rlabel metal2 s 349222 -960 349334 480 4 la_data_in[63]
port 231 nsew
rlabel metal2 s 352810 -960 352922 480 4 la_data_in[64]
port 232 nsew
rlabel metal2 s 356306 -960 356418 480 4 la_data_in[65]
port 233 nsew
rlabel metal2 s 359894 -960 360006 480 4 la_data_in[66]
port 234 nsew
rlabel metal2 s 363482 -960 363594 480 4 la_data_in[67]
port 235 nsew
rlabel metal2 s 366978 -960 367090 480 4 la_data_in[68]
port 236 nsew
rlabel metal2 s 370566 -960 370678 480 4 la_data_in[69]
port 237 nsew
rlabel metal2 s 147098 -960 147210 480 4 la_data_in[6]
port 238 nsew
rlabel metal2 s 374062 -960 374174 480 4 la_data_in[70]
port 239 nsew
rlabel metal2 s 377650 -960 377762 480 4 la_data_in[71]
port 240 nsew
rlabel metal2 s 381146 -960 381258 480 4 la_data_in[72]
port 241 nsew
rlabel metal2 s 384734 -960 384846 480 4 la_data_in[73]
port 242 nsew
rlabel metal2 s 388230 -960 388342 480 4 la_data_in[74]
port 243 nsew
rlabel metal2 s 391818 -960 391930 480 4 la_data_in[75]
port 244 nsew
rlabel metal2 s 395314 -960 395426 480 4 la_data_in[76]
port 245 nsew
rlabel metal2 s 398902 -960 399014 480 4 la_data_in[77]
port 246 nsew
rlabel metal2 s 402490 -960 402602 480 4 la_data_in[78]
port 247 nsew
rlabel metal2 s 405986 -960 406098 480 4 la_data_in[79]
port 248 nsew
rlabel metal2 s 150594 -960 150706 480 4 la_data_in[7]
port 249 nsew
rlabel metal2 s 409574 -960 409686 480 4 la_data_in[80]
port 250 nsew
rlabel metal2 s 413070 -960 413182 480 4 la_data_in[81]
port 251 nsew
rlabel metal2 s 416658 -960 416770 480 4 la_data_in[82]
port 252 nsew
rlabel metal2 s 420154 -960 420266 480 4 la_data_in[83]
port 253 nsew
rlabel metal2 s 423742 -960 423854 480 4 la_data_in[84]
port 254 nsew
rlabel metal2 s 427238 -960 427350 480 4 la_data_in[85]
port 255 nsew
rlabel metal2 s 430826 -960 430938 480 4 la_data_in[86]
port 256 nsew
rlabel metal2 s 434414 -960 434526 480 4 la_data_in[87]
port 257 nsew
rlabel metal2 s 437910 -960 438022 480 4 la_data_in[88]
port 258 nsew
rlabel metal2 s 441498 -960 441610 480 4 la_data_in[89]
port 259 nsew
rlabel metal2 s 154182 -960 154294 480 4 la_data_in[8]
port 260 nsew
rlabel metal2 s 444994 -960 445106 480 4 la_data_in[90]
port 261 nsew
rlabel metal2 s 448582 -960 448694 480 4 la_data_in[91]
port 262 nsew
rlabel metal2 s 452078 -960 452190 480 4 la_data_in[92]
port 263 nsew
rlabel metal2 s 455666 -960 455778 480 4 la_data_in[93]
port 264 nsew
rlabel metal2 s 459162 -960 459274 480 4 la_data_in[94]
port 265 nsew
rlabel metal2 s 462750 -960 462862 480 4 la_data_in[95]
port 266 nsew
rlabel metal2 s 466246 -960 466358 480 4 la_data_in[96]
port 267 nsew
rlabel metal2 s 469834 -960 469946 480 4 la_data_in[97]
port 268 nsew
rlabel metal2 s 473422 -960 473534 480 4 la_data_in[98]
port 269 nsew
rlabel metal2 s 476918 -960 477030 480 4 la_data_in[99]
port 270 nsew
rlabel metal2 s 157770 -960 157882 480 4 la_data_in[9]
port 271 nsew
rlabel metal2 s 126950 -960 127062 480 4 la_data_out[0]
port 272 nsew
rlabel metal2 s 481702 -960 481814 480 4 la_data_out[100]
port 273 nsew
rlabel metal2 s 485198 -960 485310 480 4 la_data_out[101]
port 274 nsew
rlabel metal2 s 488786 -960 488898 480 4 la_data_out[102]
port 275 nsew
rlabel metal2 s 492282 -960 492394 480 4 la_data_out[103]
port 276 nsew
rlabel metal2 s 495870 -960 495982 480 4 la_data_out[104]
port 277 nsew
rlabel metal2 s 499366 -960 499478 480 4 la_data_out[105]
port 278 nsew
rlabel metal2 s 502954 -960 503066 480 4 la_data_out[106]
port 279 nsew
rlabel metal2 s 506450 -960 506562 480 4 la_data_out[107]
port 280 nsew
rlabel metal2 s 510038 -960 510150 480 4 la_data_out[108]
port 281 nsew
rlabel metal2 s 513534 -960 513646 480 4 la_data_out[109]
port 282 nsew
rlabel metal2 s 162462 -960 162574 480 4 la_data_out[10]
port 283 nsew
rlabel metal2 s 517122 -960 517234 480 4 la_data_out[110]
port 284 nsew
rlabel metal2 s 520710 -960 520822 480 4 la_data_out[111]
port 285 nsew
rlabel metal2 s 524206 -960 524318 480 4 la_data_out[112]
port 286 nsew
rlabel metal2 s 527794 -960 527906 480 4 la_data_out[113]
port 287 nsew
rlabel metal2 s 531290 -960 531402 480 4 la_data_out[114]
port 288 nsew
rlabel metal2 s 534878 -960 534990 480 4 la_data_out[115]
port 289 nsew
rlabel metal2 s 538374 -960 538486 480 4 la_data_out[116]
port 290 nsew
rlabel metal2 s 541962 -960 542074 480 4 la_data_out[117]
port 291 nsew
rlabel metal2 s 545458 -960 545570 480 4 la_data_out[118]
port 292 nsew
rlabel metal2 s 549046 -960 549158 480 4 la_data_out[119]
port 293 nsew
rlabel metal2 s 166050 -960 166162 480 4 la_data_out[11]
port 294 nsew
rlabel metal2 s 552634 -960 552746 480 4 la_data_out[120]
port 295 nsew
rlabel metal2 s 556130 -960 556242 480 4 la_data_out[121]
port 296 nsew
rlabel metal2 s 559718 -960 559830 480 4 la_data_out[122]
port 297 nsew
rlabel metal2 s 563214 -960 563326 480 4 la_data_out[123]
port 298 nsew
rlabel metal2 s 566802 -960 566914 480 4 la_data_out[124]
port 299 nsew
rlabel metal2 s 570298 -960 570410 480 4 la_data_out[125]
port 300 nsew
rlabel metal2 s 573886 -960 573998 480 4 la_data_out[126]
port 301 nsew
rlabel metal2 s 577382 -960 577494 480 4 la_data_out[127]
port 302 nsew
rlabel metal2 s 169546 -960 169658 480 4 la_data_out[12]
port 303 nsew
rlabel metal2 s 173134 -960 173246 480 4 la_data_out[13]
port 304 nsew
rlabel metal2 s 176630 -960 176742 480 4 la_data_out[14]
port 305 nsew
rlabel metal2 s 180218 -960 180330 480 4 la_data_out[15]
port 306 nsew
rlabel metal2 s 183714 -960 183826 480 4 la_data_out[16]
port 307 nsew
rlabel metal2 s 187302 -960 187414 480 4 la_data_out[17]
port 308 nsew
rlabel metal2 s 190798 -960 190910 480 4 la_data_out[18]
port 309 nsew
rlabel metal2 s 194386 -960 194498 480 4 la_data_out[19]
port 310 nsew
rlabel metal2 s 130538 -960 130650 480 4 la_data_out[1]
port 311 nsew
rlabel metal2 s 197882 -960 197994 480 4 la_data_out[20]
port 312 nsew
rlabel metal2 s 201470 -960 201582 480 4 la_data_out[21]
port 313 nsew
rlabel metal2 s 205058 -960 205170 480 4 la_data_out[22]
port 314 nsew
rlabel metal2 s 208554 -960 208666 480 4 la_data_out[23]
port 315 nsew
rlabel metal2 s 212142 -960 212254 480 4 la_data_out[24]
port 316 nsew
rlabel metal2 s 215638 -960 215750 480 4 la_data_out[25]
port 317 nsew
rlabel metal2 s 219226 -960 219338 480 4 la_data_out[26]
port 318 nsew
rlabel metal2 s 222722 -960 222834 480 4 la_data_out[27]
port 319 nsew
rlabel metal2 s 226310 -960 226422 480 4 la_data_out[28]
port 320 nsew
rlabel metal2 s 229806 -960 229918 480 4 la_data_out[29]
port 321 nsew
rlabel metal2 s 134126 -960 134238 480 4 la_data_out[2]
port 322 nsew
rlabel metal2 s 233394 -960 233506 480 4 la_data_out[30]
port 323 nsew
rlabel metal2 s 236982 -960 237094 480 4 la_data_out[31]
port 324 nsew
rlabel metal2 s 240478 -960 240590 480 4 la_data_out[32]
port 325 nsew
rlabel metal2 s 244066 -960 244178 480 4 la_data_out[33]
port 326 nsew
rlabel metal2 s 247562 -960 247674 480 4 la_data_out[34]
port 327 nsew
rlabel metal2 s 251150 -960 251262 480 4 la_data_out[35]
port 328 nsew
rlabel metal2 s 254646 -960 254758 480 4 la_data_out[36]
port 329 nsew
rlabel metal2 s 258234 -960 258346 480 4 la_data_out[37]
port 330 nsew
rlabel metal2 s 261730 -960 261842 480 4 la_data_out[38]
port 331 nsew
rlabel metal2 s 265318 -960 265430 480 4 la_data_out[39]
port 332 nsew
rlabel metal2 s 137622 -960 137734 480 4 la_data_out[3]
port 333 nsew
rlabel metal2 s 268814 -960 268926 480 4 la_data_out[40]
port 334 nsew
rlabel metal2 s 272402 -960 272514 480 4 la_data_out[41]
port 335 nsew
rlabel metal2 s 275990 -960 276102 480 4 la_data_out[42]
port 336 nsew
rlabel metal2 s 279486 -960 279598 480 4 la_data_out[43]
port 337 nsew
rlabel metal2 s 283074 -960 283186 480 4 la_data_out[44]
port 338 nsew
rlabel metal2 s 286570 -960 286682 480 4 la_data_out[45]
port 339 nsew
rlabel metal2 s 290158 -960 290270 480 4 la_data_out[46]
port 340 nsew
rlabel metal2 s 293654 -960 293766 480 4 la_data_out[47]
port 341 nsew
rlabel metal2 s 297242 -960 297354 480 4 la_data_out[48]
port 342 nsew
rlabel metal2 s 300738 -960 300850 480 4 la_data_out[49]
port 343 nsew
rlabel metal2 s 141210 -960 141322 480 4 la_data_out[4]
port 344 nsew
rlabel metal2 s 304326 -960 304438 480 4 la_data_out[50]
port 345 nsew
rlabel metal2 s 307914 -960 308026 480 4 la_data_out[51]
port 346 nsew
rlabel metal2 s 311410 -960 311522 480 4 la_data_out[52]
port 347 nsew
rlabel metal2 s 314998 -960 315110 480 4 la_data_out[53]
port 348 nsew
rlabel metal2 s 318494 -960 318606 480 4 la_data_out[54]
port 349 nsew
rlabel metal2 s 322082 -960 322194 480 4 la_data_out[55]
port 350 nsew
rlabel metal2 s 325578 -960 325690 480 4 la_data_out[56]
port 351 nsew
rlabel metal2 s 329166 -960 329278 480 4 la_data_out[57]
port 352 nsew
rlabel metal2 s 332662 -960 332774 480 4 la_data_out[58]
port 353 nsew
rlabel metal2 s 336250 -960 336362 480 4 la_data_out[59]
port 354 nsew
rlabel metal2 s 144706 -960 144818 480 4 la_data_out[5]
port 355 nsew
rlabel metal2 s 339838 -960 339950 480 4 la_data_out[60]
port 356 nsew
rlabel metal2 s 343334 -960 343446 480 4 la_data_out[61]
port 357 nsew
rlabel metal2 s 346922 -960 347034 480 4 la_data_out[62]
port 358 nsew
rlabel metal2 s 350418 -960 350530 480 4 la_data_out[63]
port 359 nsew
rlabel metal2 s 354006 -960 354118 480 4 la_data_out[64]
port 360 nsew
rlabel metal2 s 357502 -960 357614 480 4 la_data_out[65]
port 361 nsew
rlabel metal2 s 361090 -960 361202 480 4 la_data_out[66]
port 362 nsew
rlabel metal2 s 364586 -960 364698 480 4 la_data_out[67]
port 363 nsew
rlabel metal2 s 368174 -960 368286 480 4 la_data_out[68]
port 364 nsew
rlabel metal2 s 371670 -960 371782 480 4 la_data_out[69]
port 365 nsew
rlabel metal2 s 148294 -960 148406 480 4 la_data_out[6]
port 366 nsew
rlabel metal2 s 375258 -960 375370 480 4 la_data_out[70]
port 367 nsew
rlabel metal2 s 378846 -960 378958 480 4 la_data_out[71]
port 368 nsew
rlabel metal2 s 382342 -960 382454 480 4 la_data_out[72]
port 369 nsew
rlabel metal2 s 385930 -960 386042 480 4 la_data_out[73]
port 370 nsew
rlabel metal2 s 389426 -960 389538 480 4 la_data_out[74]
port 371 nsew
rlabel metal2 s 393014 -960 393126 480 4 la_data_out[75]
port 372 nsew
rlabel metal2 s 396510 -960 396622 480 4 la_data_out[76]
port 373 nsew
rlabel metal2 s 400098 -960 400210 480 4 la_data_out[77]
port 374 nsew
rlabel metal2 s 403594 -960 403706 480 4 la_data_out[78]
port 375 nsew
rlabel metal2 s 407182 -960 407294 480 4 la_data_out[79]
port 376 nsew
rlabel metal2 s 151790 -960 151902 480 4 la_data_out[7]
port 377 nsew
rlabel metal2 s 410770 -960 410882 480 4 la_data_out[80]
port 378 nsew
rlabel metal2 s 414266 -960 414378 480 4 la_data_out[81]
port 379 nsew
rlabel metal2 s 417854 -960 417966 480 4 la_data_out[82]
port 380 nsew
rlabel metal2 s 421350 -960 421462 480 4 la_data_out[83]
port 381 nsew
rlabel metal2 s 424938 -960 425050 480 4 la_data_out[84]
port 382 nsew
rlabel metal2 s 428434 -960 428546 480 4 la_data_out[85]
port 383 nsew
rlabel metal2 s 432022 -960 432134 480 4 la_data_out[86]
port 384 nsew
rlabel metal2 s 435518 -960 435630 480 4 la_data_out[87]
port 385 nsew
rlabel metal2 s 439106 -960 439218 480 4 la_data_out[88]
port 386 nsew
rlabel metal2 s 442602 -960 442714 480 4 la_data_out[89]
port 387 nsew
rlabel metal2 s 155378 -960 155490 480 4 la_data_out[8]
port 388 nsew
rlabel metal2 s 446190 -960 446302 480 4 la_data_out[90]
port 389 nsew
rlabel metal2 s 449778 -960 449890 480 4 la_data_out[91]
port 390 nsew
rlabel metal2 s 453274 -960 453386 480 4 la_data_out[92]
port 391 nsew
rlabel metal2 s 456862 -960 456974 480 4 la_data_out[93]
port 392 nsew
rlabel metal2 s 460358 -960 460470 480 4 la_data_out[94]
port 393 nsew
rlabel metal2 s 463946 -960 464058 480 4 la_data_out[95]
port 394 nsew
rlabel metal2 s 467442 -960 467554 480 4 la_data_out[96]
port 395 nsew
rlabel metal2 s 471030 -960 471142 480 4 la_data_out[97]
port 396 nsew
rlabel metal2 s 474526 -960 474638 480 4 la_data_out[98]
port 397 nsew
rlabel metal2 s 478114 -960 478226 480 4 la_data_out[99]
port 398 nsew
rlabel metal2 s 158874 -960 158986 480 4 la_data_out[9]
port 399 nsew
rlabel metal2 s 128146 -960 128258 480 4 la_oenb[0]
port 400 nsew
rlabel metal2 s 482806 -960 482918 480 4 la_oenb[100]
port 401 nsew
rlabel metal2 s 486394 -960 486506 480 4 la_oenb[101]
port 402 nsew
rlabel metal2 s 489890 -960 490002 480 4 la_oenb[102]
port 403 nsew
rlabel metal2 s 493478 -960 493590 480 4 la_oenb[103]
port 404 nsew
rlabel metal2 s 497066 -960 497178 480 4 la_oenb[104]
port 405 nsew
rlabel metal2 s 500562 -960 500674 480 4 la_oenb[105]
port 406 nsew
rlabel metal2 s 504150 -960 504262 480 4 la_oenb[106]
port 407 nsew
rlabel metal2 s 507646 -960 507758 480 4 la_oenb[107]
port 408 nsew
rlabel metal2 s 511234 -960 511346 480 4 la_oenb[108]
port 409 nsew
rlabel metal2 s 514730 -960 514842 480 4 la_oenb[109]
port 410 nsew
rlabel metal2 s 163658 -960 163770 480 4 la_oenb[10]
port 411 nsew
rlabel metal2 s 518318 -960 518430 480 4 la_oenb[110]
port 412 nsew
rlabel metal2 s 521814 -960 521926 480 4 la_oenb[111]
port 413 nsew
rlabel metal2 s 525402 -960 525514 480 4 la_oenb[112]
port 414 nsew
rlabel metal2 s 528990 -960 529102 480 4 la_oenb[113]
port 415 nsew
rlabel metal2 s 532486 -960 532598 480 4 la_oenb[114]
port 416 nsew
rlabel metal2 s 536074 -960 536186 480 4 la_oenb[115]
port 417 nsew
rlabel metal2 s 539570 -960 539682 480 4 la_oenb[116]
port 418 nsew
rlabel metal2 s 543158 -960 543270 480 4 la_oenb[117]
port 419 nsew
rlabel metal2 s 546654 -960 546766 480 4 la_oenb[118]
port 420 nsew
rlabel metal2 s 550242 -960 550354 480 4 la_oenb[119]
port 421 nsew
rlabel metal2 s 167154 -960 167266 480 4 la_oenb[11]
port 422 nsew
rlabel metal2 s 553738 -960 553850 480 4 la_oenb[120]
port 423 nsew
rlabel metal2 s 557326 -960 557438 480 4 la_oenb[121]
port 424 nsew
rlabel metal2 s 560822 -960 560934 480 4 la_oenb[122]
port 425 nsew
rlabel metal2 s 564410 -960 564522 480 4 la_oenb[123]
port 426 nsew
rlabel metal2 s 567998 -960 568110 480 4 la_oenb[124]
port 427 nsew
rlabel metal2 s 571494 -960 571606 480 4 la_oenb[125]
port 428 nsew
rlabel metal2 s 575082 -960 575194 480 4 la_oenb[126]
port 429 nsew
rlabel metal2 s 578578 -960 578690 480 4 la_oenb[127]
port 430 nsew
rlabel metal2 s 170742 -960 170854 480 4 la_oenb[12]
port 431 nsew
rlabel metal2 s 174238 -960 174350 480 4 la_oenb[13]
port 432 nsew
rlabel metal2 s 177826 -960 177938 480 4 la_oenb[14]
port 433 nsew
rlabel metal2 s 181414 -960 181526 480 4 la_oenb[15]
port 434 nsew
rlabel metal2 s 184910 -960 185022 480 4 la_oenb[16]
port 435 nsew
rlabel metal2 s 188498 -960 188610 480 4 la_oenb[17]
port 436 nsew
rlabel metal2 s 191994 -960 192106 480 4 la_oenb[18]
port 437 nsew
rlabel metal2 s 195582 -960 195694 480 4 la_oenb[19]
port 438 nsew
rlabel metal2 s 131734 -960 131846 480 4 la_oenb[1]
port 439 nsew
rlabel metal2 s 199078 -960 199190 480 4 la_oenb[20]
port 440 nsew
rlabel metal2 s 202666 -960 202778 480 4 la_oenb[21]
port 441 nsew
rlabel metal2 s 206162 -960 206274 480 4 la_oenb[22]
port 442 nsew
rlabel metal2 s 209750 -960 209862 480 4 la_oenb[23]
port 443 nsew
rlabel metal2 s 213338 -960 213450 480 4 la_oenb[24]
port 444 nsew
rlabel metal2 s 216834 -960 216946 480 4 la_oenb[25]
port 445 nsew
rlabel metal2 s 220422 -960 220534 480 4 la_oenb[26]
port 446 nsew
rlabel metal2 s 223918 -960 224030 480 4 la_oenb[27]
port 447 nsew
rlabel metal2 s 227506 -960 227618 480 4 la_oenb[28]
port 448 nsew
rlabel metal2 s 231002 -960 231114 480 4 la_oenb[29]
port 449 nsew
rlabel metal2 s 135230 -960 135342 480 4 la_oenb[2]
port 450 nsew
rlabel metal2 s 234590 -960 234702 480 4 la_oenb[30]
port 451 nsew
rlabel metal2 s 238086 -960 238198 480 4 la_oenb[31]
port 452 nsew
rlabel metal2 s 241674 -960 241786 480 4 la_oenb[32]
port 453 nsew
rlabel metal2 s 245170 -960 245282 480 4 la_oenb[33]
port 454 nsew
rlabel metal2 s 248758 -960 248870 480 4 la_oenb[34]
port 455 nsew
rlabel metal2 s 252346 -960 252458 480 4 la_oenb[35]
port 456 nsew
rlabel metal2 s 255842 -960 255954 480 4 la_oenb[36]
port 457 nsew
rlabel metal2 s 259430 -960 259542 480 4 la_oenb[37]
port 458 nsew
rlabel metal2 s 262926 -960 263038 480 4 la_oenb[38]
port 459 nsew
rlabel metal2 s 266514 -960 266626 480 4 la_oenb[39]
port 460 nsew
rlabel metal2 s 138818 -960 138930 480 4 la_oenb[3]
port 461 nsew
rlabel metal2 s 270010 -960 270122 480 4 la_oenb[40]
port 462 nsew
rlabel metal2 s 273598 -960 273710 480 4 la_oenb[41]
port 463 nsew
rlabel metal2 s 277094 -960 277206 480 4 la_oenb[42]
port 464 nsew
rlabel metal2 s 280682 -960 280794 480 4 la_oenb[43]
port 465 nsew
rlabel metal2 s 284270 -960 284382 480 4 la_oenb[44]
port 466 nsew
rlabel metal2 s 287766 -960 287878 480 4 la_oenb[45]
port 467 nsew
rlabel metal2 s 291354 -960 291466 480 4 la_oenb[46]
port 468 nsew
rlabel metal2 s 294850 -960 294962 480 4 la_oenb[47]
port 469 nsew
rlabel metal2 s 298438 -960 298550 480 4 la_oenb[48]
port 470 nsew
rlabel metal2 s 301934 -960 302046 480 4 la_oenb[49]
port 471 nsew
rlabel metal2 s 142406 -960 142518 480 4 la_oenb[4]
port 472 nsew
rlabel metal2 s 305522 -960 305634 480 4 la_oenb[50]
port 473 nsew
rlabel metal2 s 309018 -960 309130 480 4 la_oenb[51]
port 474 nsew
rlabel metal2 s 312606 -960 312718 480 4 la_oenb[52]
port 475 nsew
rlabel metal2 s 316194 -960 316306 480 4 la_oenb[53]
port 476 nsew
rlabel metal2 s 319690 -960 319802 480 4 la_oenb[54]
port 477 nsew
rlabel metal2 s 323278 -960 323390 480 4 la_oenb[55]
port 478 nsew
rlabel metal2 s 326774 -960 326886 480 4 la_oenb[56]
port 479 nsew
rlabel metal2 s 330362 -960 330474 480 4 la_oenb[57]
port 480 nsew
rlabel metal2 s 333858 -960 333970 480 4 la_oenb[58]
port 481 nsew
rlabel metal2 s 337446 -960 337558 480 4 la_oenb[59]
port 482 nsew
rlabel metal2 s 145902 -960 146014 480 4 la_oenb[5]
port 483 nsew
rlabel metal2 s 340942 -960 341054 480 4 la_oenb[60]
port 484 nsew
rlabel metal2 s 344530 -960 344642 480 4 la_oenb[61]
port 485 nsew
rlabel metal2 s 348026 -960 348138 480 4 la_oenb[62]
port 486 nsew
rlabel metal2 s 351614 -960 351726 480 4 la_oenb[63]
port 487 nsew
rlabel metal2 s 355202 -960 355314 480 4 la_oenb[64]
port 488 nsew
rlabel metal2 s 358698 -960 358810 480 4 la_oenb[65]
port 489 nsew
rlabel metal2 s 362286 -960 362398 480 4 la_oenb[66]
port 490 nsew
rlabel metal2 s 365782 -960 365894 480 4 la_oenb[67]
port 491 nsew
rlabel metal2 s 369370 -960 369482 480 4 la_oenb[68]
port 492 nsew
rlabel metal2 s 372866 -960 372978 480 4 la_oenb[69]
port 493 nsew
rlabel metal2 s 149490 -960 149602 480 4 la_oenb[6]
port 494 nsew
rlabel metal2 s 376454 -960 376566 480 4 la_oenb[70]
port 495 nsew
rlabel metal2 s 379950 -960 380062 480 4 la_oenb[71]
port 496 nsew
rlabel metal2 s 383538 -960 383650 480 4 la_oenb[72]
port 497 nsew
rlabel metal2 s 387126 -960 387238 480 4 la_oenb[73]
port 498 nsew
rlabel metal2 s 390622 -960 390734 480 4 la_oenb[74]
port 499 nsew
rlabel metal2 s 394210 -960 394322 480 4 la_oenb[75]
port 500 nsew
rlabel metal2 s 397706 -960 397818 480 4 la_oenb[76]
port 501 nsew
rlabel metal2 s 401294 -960 401406 480 4 la_oenb[77]
port 502 nsew
rlabel metal2 s 404790 -960 404902 480 4 la_oenb[78]
port 503 nsew
rlabel metal2 s 408378 -960 408490 480 4 la_oenb[79]
port 504 nsew
rlabel metal2 s 152986 -960 153098 480 4 la_oenb[7]
port 505 nsew
rlabel metal2 s 411874 -960 411986 480 4 la_oenb[80]
port 506 nsew
rlabel metal2 s 415462 -960 415574 480 4 la_oenb[81]
port 507 nsew
rlabel metal2 s 418958 -960 419070 480 4 la_oenb[82]
port 508 nsew
rlabel metal2 s 422546 -960 422658 480 4 la_oenb[83]
port 509 nsew
rlabel metal2 s 426134 -960 426246 480 4 la_oenb[84]
port 510 nsew
rlabel metal2 s 429630 -960 429742 480 4 la_oenb[85]
port 511 nsew
rlabel metal2 s 433218 -960 433330 480 4 la_oenb[86]
port 512 nsew
rlabel metal2 s 436714 -960 436826 480 4 la_oenb[87]
port 513 nsew
rlabel metal2 s 440302 -960 440414 480 4 la_oenb[88]
port 514 nsew
rlabel metal2 s 443798 -960 443910 480 4 la_oenb[89]
port 515 nsew
rlabel metal2 s 156574 -960 156686 480 4 la_oenb[8]
port 516 nsew
rlabel metal2 s 447386 -960 447498 480 4 la_oenb[90]
port 517 nsew
rlabel metal2 s 450882 -960 450994 480 4 la_oenb[91]
port 518 nsew
rlabel metal2 s 454470 -960 454582 480 4 la_oenb[92]
port 519 nsew
rlabel metal2 s 458058 -960 458170 480 4 la_oenb[93]
port 520 nsew
rlabel metal2 s 461554 -960 461666 480 4 la_oenb[94]
port 521 nsew
rlabel metal2 s 465142 -960 465254 480 4 la_oenb[95]
port 522 nsew
rlabel metal2 s 468638 -960 468750 480 4 la_oenb[96]
port 523 nsew
rlabel metal2 s 472226 -960 472338 480 4 la_oenb[97]
port 524 nsew
rlabel metal2 s 475722 -960 475834 480 4 la_oenb[98]
port 525 nsew
rlabel metal2 s 479310 -960 479422 480 4 la_oenb[99]
port 526 nsew
rlabel metal2 s 160070 -960 160182 480 4 la_oenb[9]
port 527 nsew
rlabel metal2 s 579774 -960 579886 480 4 user_clock2
port 528 nsew
rlabel metal2 s 580970 -960 581082 480 4 user_irq[0]
port 529 nsew
rlabel metal2 s 582166 -960 582278 480 4 user_irq[1]
port 530 nsew
rlabel metal2 s 583362 -960 583474 480 4 user_irq[2]
port 531 nsew
rlabel metal5 s -2006 -934 585930 -314 4 vccd1
port 532 nsew
rlabel metal5 s -2966 2866 586890 3486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 38866 586890 39486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 74866 586890 75486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 110866 586890 111486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 146866 586890 147486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 182866 586890 183486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 218866 586890 219486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 254866 586890 255486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 290866 586890 291486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 326866 586890 327486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 362866 586890 363486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 398866 586890 399486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 434866 586890 435486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 470866 586890 471486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 506866 586890 507486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 542866 586890 543486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 578866 586890 579486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 614866 586890 615486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 650866 586890 651486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 686866 586890 687486 4 vccd1
port 532 nsew
rlabel metal5 s -2006 704250 585930 704870 4 vccd1
port 532 nsew
rlabel metal4 s 253794 -1894 254414 338000 4 vccd1
port 532 nsew
rlabel metal4 s 289794 -1894 290414 338000 4 vccd1
port 532 nsew
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 532 nsew
rlabel metal4 s 585310 -934 585930 704870 4 vccd1
port 532 nsew
rlabel metal4 s 1794 -1894 2414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 37794 -1894 38414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 73794 -1894 74414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 109794 -1894 110414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 145794 -1894 146414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 181794 -1894 182414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 217794 -1894 218414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 253794 378000 254414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 289794 378000 290414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 325794 -1894 326414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 361794 -1894 362414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 397794 -1894 398414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 433794 -1894 434414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 469794 -1894 470414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 505794 -1894 506414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 541794 -1894 542414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 577794 -1894 578414 705830 4 vccd1
port 532 nsew
rlabel metal5 s -3926 -2854 587850 -2234 4 vccd2
port 533 nsew
rlabel metal5 s -4886 6586 588810 7206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 42586 588810 43206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 78586 588810 79206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 114586 588810 115206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 150586 588810 151206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 186586 588810 187206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 222586 588810 223206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 258586 588810 259206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 294586 588810 295206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 330586 588810 331206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 366586 588810 367206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 402586 588810 403206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 438586 588810 439206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 474586 588810 475206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 510586 588810 511206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 546586 588810 547206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 582586 588810 583206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 618586 588810 619206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 654586 588810 655206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 690586 588810 691206 4 vccd2
port 533 nsew
rlabel metal5 s -3926 706170 587850 706790 4 vccd2
port 533 nsew
rlabel metal4 s 257514 -3814 258134 336000 4 vccd2
port 533 nsew
rlabel metal4 s 293514 -3814 294134 336000 4 vccd2
port 533 nsew
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 533 nsew
rlabel metal4 s 587230 -2854 587850 706790 4 vccd2
port 533 nsew
rlabel metal4 s 5514 -3814 6134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 41514 -3814 42134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 77514 -3814 78134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 113514 -3814 114134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 149514 -3814 150134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 185514 -3814 186134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 221514 -3814 222134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 257514 380000 258134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 293514 380000 294134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 329514 -3814 330134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 365514 -3814 366134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 401514 -3814 402134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 437514 -3814 438134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 473514 -3814 474134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 509514 -3814 510134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 545514 -3814 546134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 581514 -3814 582134 707750 4 vccd2
port 533 nsew
rlabel metal5 s -5846 -4774 589770 -4154 4 vdda1
port 534 nsew
rlabel metal5 s -6806 10306 590730 10926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 46306 590730 46926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 82306 590730 82926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 118306 590730 118926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 154306 590730 154926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 190306 590730 190926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 226306 590730 226926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 262306 590730 262926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 298306 590730 298926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 334306 590730 334926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 370306 590730 370926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 406306 590730 406926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 442306 590730 442926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 478306 590730 478926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 514306 590730 514926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 550306 590730 550926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 586306 590730 586926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 622306 590730 622926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 658306 590730 658926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 694306 590730 694926 4 vdda1
port 534 nsew
rlabel metal5 s -5846 708090 589770 708710 4 vdda1
port 534 nsew
rlabel metal4 s 261234 -5734 261854 336000 4 vdda1
port 534 nsew
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 534 nsew
rlabel metal4 s 589150 -4774 589770 708710 4 vdda1
port 534 nsew
rlabel metal4 s 9234 -5734 9854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 45234 -5734 45854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 81234 -5734 81854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 117234 -5734 117854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 153234 -5734 153854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 189234 -5734 189854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 225234 -5734 225854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 261234 380000 261854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 297234 -5734 297854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 333234 -5734 333854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 369234 -5734 369854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 405234 -5734 405854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 441234 -5734 441854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 477234 -5734 477854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 513234 -5734 513854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 549234 -5734 549854 709670 4 vdda1
port 534 nsew
rlabel metal5 s -7766 -6694 591690 -6074 4 vdda2
port 535 nsew
rlabel metal5 s -8726 14026 592650 14646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 50026 592650 50646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 86026 592650 86646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 122026 592650 122646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 158026 592650 158646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 194026 592650 194646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 230026 592650 230646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 266026 592650 266646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 302026 592650 302646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 338026 592650 338646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 374026 592650 374646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 410026 592650 410646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 446026 592650 446646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 482026 592650 482646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 518026 592650 518646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 554026 592650 554646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 590026 592650 590646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 626026 592650 626646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 662026 592650 662646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 698026 592650 698646 4 vdda2
port 535 nsew
rlabel metal5 s -7766 710010 591690 710630 4 vdda2
port 535 nsew
rlabel metal4 s 264954 -7654 265574 336000 4 vdda2
port 535 nsew
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 535 nsew
rlabel metal4 s 591070 -6694 591690 710630 4 vdda2
port 535 nsew
rlabel metal4 s 12954 -7654 13574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 48954 -7654 49574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 84954 -7654 85574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 120954 -7654 121574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 156954 -7654 157574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 192954 -7654 193574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 228954 -7654 229574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 264954 380000 265574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 300954 -7654 301574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 336954 -7654 337574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 372954 -7654 373574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 408954 -7654 409574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 444954 -7654 445574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 480954 -7654 481574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 516954 -7654 517574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 552954 -7654 553574 711590 4 vdda2
port 535 nsew
rlabel metal5 s -6806 -5734 590730 -5114 4 vssa1
port 536 nsew
rlabel metal5 s -6806 28306 590730 28926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 64306 590730 64926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 100306 590730 100926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 136306 590730 136926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 172306 590730 172926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 208306 590730 208926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 244306 590730 244926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 280306 590730 280926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 316306 590730 316926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 352306 590730 352926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 388306 590730 388926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 424306 590730 424926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 460306 590730 460926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 496306 590730 496926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 532306 590730 532926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 568306 590730 568926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 604306 590730 604926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 640306 590730 640926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 676306 590730 676926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 709050 590730 709670 4 vssa1
port 536 nsew
rlabel metal4 s 243234 -5734 243854 336000 4 vssa1
port 536 nsew
rlabel metal4 s 279234 -5734 279854 336000 4 vssa1
port 536 nsew
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 536 nsew
rlabel metal4 s 27234 -5734 27854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 63234 -5734 63854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 99234 -5734 99854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 135234 -5734 135854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 171234 -5734 171854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 207234 -5734 207854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 243234 380000 243854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 279234 380000 279854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 315234 -5734 315854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 351234 -5734 351854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 387234 -5734 387854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 423234 -5734 423854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 459234 -5734 459854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 495234 -5734 495854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 531234 -5734 531854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 567234 -5734 567854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 590110 -5734 590730 709670 4 vssa1
port 536 nsew
rlabel metal5 s -8726 -7654 592650 -7034 4 vssa2
port 537 nsew
rlabel metal5 s -8726 32026 592650 32646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 68026 592650 68646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 104026 592650 104646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 140026 592650 140646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 176026 592650 176646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 212026 592650 212646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 248026 592650 248646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 284026 592650 284646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 320026 592650 320646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 356026 592650 356646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 392026 592650 392646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 428026 592650 428646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 464026 592650 464646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 500026 592650 500646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 536026 592650 536646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 572026 592650 572646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 608026 592650 608646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 644026 592650 644646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 680026 592650 680646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 710970 592650 711590 4 vssa2
port 537 nsew
rlabel metal4 s 246954 -7654 247574 336000 4 vssa2
port 537 nsew
rlabel metal4 s 282954 -7654 283574 336000 4 vssa2
port 537 nsew
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 537 nsew
rlabel metal4 s 30954 -7654 31574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 66954 -7654 67574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 102954 -7654 103574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 138954 -7654 139574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 174954 -7654 175574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 210954 -7654 211574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 246954 380000 247574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 282954 380000 283574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 318954 -7654 319574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 354954 -7654 355574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 390954 -7654 391574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 426954 -7654 427574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 462954 -7654 463574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 498954 -7654 499574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 534954 -7654 535574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 570954 -7654 571574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 592030 -7654 592650 711590 4 vssa2
port 537 nsew
rlabel metal5 s -2966 -1894 586890 -1274 4 vssd1
port 538 nsew
rlabel metal5 s -2966 20866 586890 21486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 56866 586890 57486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 92866 586890 93486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 128866 586890 129486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 164866 586890 165486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 200866 586890 201486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 236866 586890 237486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 272866 586890 273486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 308866 586890 309486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 344866 586890 345486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 380866 586890 381486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 416866 586890 417486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 452866 586890 453486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 488866 586890 489486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 524866 586890 525486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 560866 586890 561486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 596866 586890 597486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 632866 586890 633486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 668866 586890 669486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 705210 586890 705830 4 vssd1
port 538 nsew
rlabel metal4 s 235794 -1894 236414 338000 4 vssd1
port 538 nsew
rlabel metal4 s 271794 -1894 272414 338000 4 vssd1
port 538 nsew
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 538 nsew
rlabel metal4 s 19794 -1894 20414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 55794 -1894 56414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 91794 -1894 92414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 127794 -1894 128414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 163794 -1894 164414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 199794 -1894 200414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 235794 378000 236414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 271794 378000 272414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 307794 -1894 308414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 343794 -1894 344414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 379794 -1894 380414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 415794 -1894 416414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 451794 -1894 452414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 487794 -1894 488414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 523794 -1894 524414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 559794 -1894 560414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 586270 -1894 586890 705830 4 vssd1
port 538 nsew
rlabel metal5 s -4886 -3814 588810 -3194 4 vssd2
port 539 nsew
rlabel metal5 s -4886 24586 588810 25206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 60586 588810 61206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 96586 588810 97206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 132586 588810 133206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 168586 588810 169206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 204586 588810 205206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 240586 588810 241206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 276586 588810 277206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 312586 588810 313206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 348586 588810 349206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 384586 588810 385206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 420586 588810 421206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 456586 588810 457206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 492586 588810 493206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 528586 588810 529206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 564586 588810 565206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 600586 588810 601206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 636586 588810 637206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 672586 588810 673206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 707130 588810 707750 4 vssd2
port 539 nsew
rlabel metal4 s 239514 -3814 240134 336000 4 vssd2
port 539 nsew
rlabel metal4 s 275514 -3814 276134 336000 4 vssd2
port 539 nsew
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 539 nsew
rlabel metal4 s 23514 -3814 24134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 59514 -3814 60134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 95514 -3814 96134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 131514 -3814 132134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 167514 -3814 168134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 203514 -3814 204134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 239514 380000 240134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 275514 380000 276134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 311514 -3814 312134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 347514 -3814 348134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 383514 -3814 384134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 419514 -3814 420134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 455514 -3814 456134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 491514 -3814 492134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 527514 -3814 528134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 563514 -3814 564134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 588190 -3814 588810 707750 4 vssd2
port 539 nsew
rlabel metal2 s 542 -960 654 480 4 wb_clk_i
port 540 nsew
rlabel metal2 s 1646 -960 1758 480 4 wb_rst_i
port 541 nsew
rlabel metal2 s 2842 -960 2954 480 4 wbs_ack_o
port 542 nsew
rlabel metal2 s 7626 -960 7738 480 4 wbs_adr_i[0]
port 543 nsew
rlabel metal2 s 47830 -960 47942 480 4 wbs_adr_i[10]
port 544 nsew
rlabel metal2 s 51326 -960 51438 480 4 wbs_adr_i[11]
port 545 nsew
rlabel metal2 s 54914 -960 55026 480 4 wbs_adr_i[12]
port 546 nsew
rlabel metal2 s 58410 -960 58522 480 4 wbs_adr_i[13]
port 547 nsew
rlabel metal2 s 61998 -960 62110 480 4 wbs_adr_i[14]
port 548 nsew
rlabel metal2 s 65494 -960 65606 480 4 wbs_adr_i[15]
port 549 nsew
rlabel metal2 s 69082 -960 69194 480 4 wbs_adr_i[16]
port 550 nsew
rlabel metal2 s 72578 -960 72690 480 4 wbs_adr_i[17]
port 551 nsew
rlabel metal2 s 76166 -960 76278 480 4 wbs_adr_i[18]
port 552 nsew
rlabel metal2 s 79662 -960 79774 480 4 wbs_adr_i[19]
port 553 nsew
rlabel metal2 s 12318 -960 12430 480 4 wbs_adr_i[1]
port 554 nsew
rlabel metal2 s 83250 -960 83362 480 4 wbs_adr_i[20]
port 555 nsew
rlabel metal2 s 86838 -960 86950 480 4 wbs_adr_i[21]
port 556 nsew
rlabel metal2 s 90334 -960 90446 480 4 wbs_adr_i[22]
port 557 nsew
rlabel metal2 s 93922 -960 94034 480 4 wbs_adr_i[23]
port 558 nsew
rlabel metal2 s 97418 -960 97530 480 4 wbs_adr_i[24]
port 559 nsew
rlabel metal2 s 101006 -960 101118 480 4 wbs_adr_i[25]
port 560 nsew
rlabel metal2 s 104502 -960 104614 480 4 wbs_adr_i[26]
port 561 nsew
rlabel metal2 s 108090 -960 108202 480 4 wbs_adr_i[27]
port 562 nsew
rlabel metal2 s 111586 -960 111698 480 4 wbs_adr_i[28]
port 563 nsew
rlabel metal2 s 115174 -960 115286 480 4 wbs_adr_i[29]
port 564 nsew
rlabel metal2 s 17010 -960 17122 480 4 wbs_adr_i[2]
port 565 nsew
rlabel metal2 s 118762 -960 118874 480 4 wbs_adr_i[30]
port 566 nsew
rlabel metal2 s 122258 -960 122370 480 4 wbs_adr_i[31]
port 567 nsew
rlabel metal2 s 21794 -960 21906 480 4 wbs_adr_i[3]
port 568 nsew
rlabel metal2 s 26486 -960 26598 480 4 wbs_adr_i[4]
port 569 nsew
rlabel metal2 s 30074 -960 30186 480 4 wbs_adr_i[5]
port 570 nsew
rlabel metal2 s 33570 -960 33682 480 4 wbs_adr_i[6]
port 571 nsew
rlabel metal2 s 37158 -960 37270 480 4 wbs_adr_i[7]
port 572 nsew
rlabel metal2 s 40654 -960 40766 480 4 wbs_adr_i[8]
port 573 nsew
rlabel metal2 s 44242 -960 44354 480 4 wbs_adr_i[9]
port 574 nsew
rlabel metal2 s 4038 -960 4150 480 4 wbs_cyc_i
port 575 nsew
rlabel metal2 s 8730 -960 8842 480 4 wbs_dat_i[0]
port 576 nsew
rlabel metal2 s 48934 -960 49046 480 4 wbs_dat_i[10]
port 577 nsew
rlabel metal2 s 52522 -960 52634 480 4 wbs_dat_i[11]
port 578 nsew
rlabel metal2 s 56018 -960 56130 480 4 wbs_dat_i[12]
port 579 nsew
rlabel metal2 s 59606 -960 59718 480 4 wbs_dat_i[13]
port 580 nsew
rlabel metal2 s 63194 -960 63306 480 4 wbs_dat_i[14]
port 581 nsew
rlabel metal2 s 66690 -960 66802 480 4 wbs_dat_i[15]
port 582 nsew
rlabel metal2 s 70278 -960 70390 480 4 wbs_dat_i[16]
port 583 nsew
rlabel metal2 s 73774 -960 73886 480 4 wbs_dat_i[17]
port 584 nsew
rlabel metal2 s 77362 -960 77474 480 4 wbs_dat_i[18]
port 585 nsew
rlabel metal2 s 80858 -960 80970 480 4 wbs_dat_i[19]
port 586 nsew
rlabel metal2 s 13514 -960 13626 480 4 wbs_dat_i[1]
port 587 nsew
rlabel metal2 s 84446 -960 84558 480 4 wbs_dat_i[20]
port 588 nsew
rlabel metal2 s 87942 -960 88054 480 4 wbs_dat_i[21]
port 589 nsew
rlabel metal2 s 91530 -960 91642 480 4 wbs_dat_i[22]
port 590 nsew
rlabel metal2 s 95118 -960 95230 480 4 wbs_dat_i[23]
port 591 nsew
rlabel metal2 s 98614 -960 98726 480 4 wbs_dat_i[24]
port 592 nsew
rlabel metal2 s 102202 -960 102314 480 4 wbs_dat_i[25]
port 593 nsew
rlabel metal2 s 105698 -960 105810 480 4 wbs_dat_i[26]
port 594 nsew
rlabel metal2 s 109286 -960 109398 480 4 wbs_dat_i[27]
port 595 nsew
rlabel metal2 s 112782 -960 112894 480 4 wbs_dat_i[28]
port 596 nsew
rlabel metal2 s 116370 -960 116482 480 4 wbs_dat_i[29]
port 597 nsew
rlabel metal2 s 18206 -960 18318 480 4 wbs_dat_i[2]
port 598 nsew
rlabel metal2 s 119866 -960 119978 480 4 wbs_dat_i[30]
port 599 nsew
rlabel metal2 s 123454 -960 123566 480 4 wbs_dat_i[31]
port 600 nsew
rlabel metal2 s 22990 -960 23102 480 4 wbs_dat_i[3]
port 601 nsew
rlabel metal2 s 27682 -960 27794 480 4 wbs_dat_i[4]
port 602 nsew
rlabel metal2 s 31270 -960 31382 480 4 wbs_dat_i[5]
port 603 nsew
rlabel metal2 s 34766 -960 34878 480 4 wbs_dat_i[6]
port 604 nsew
rlabel metal2 s 38354 -960 38466 480 4 wbs_dat_i[7]
port 605 nsew
rlabel metal2 s 41850 -960 41962 480 4 wbs_dat_i[8]
port 606 nsew
rlabel metal2 s 45438 -960 45550 480 4 wbs_dat_i[9]
port 607 nsew
rlabel metal2 s 9926 -960 10038 480 4 wbs_dat_o[0]
port 608 nsew
rlabel metal2 s 50130 -960 50242 480 4 wbs_dat_o[10]
port 609 nsew
rlabel metal2 s 53718 -960 53830 480 4 wbs_dat_o[11]
port 610 nsew
rlabel metal2 s 57214 -960 57326 480 4 wbs_dat_o[12]
port 611 nsew
rlabel metal2 s 60802 -960 60914 480 4 wbs_dat_o[13]
port 612 nsew
rlabel metal2 s 64298 -960 64410 480 4 wbs_dat_o[14]
port 613 nsew
rlabel metal2 s 67886 -960 67998 480 4 wbs_dat_o[15]
port 614 nsew
rlabel metal2 s 71474 -960 71586 480 4 wbs_dat_o[16]
port 615 nsew
rlabel metal2 s 74970 -960 75082 480 4 wbs_dat_o[17]
port 616 nsew
rlabel metal2 s 78558 -960 78670 480 4 wbs_dat_o[18]
port 617 nsew
rlabel metal2 s 82054 -960 82166 480 4 wbs_dat_o[19]
port 618 nsew
rlabel metal2 s 14710 -960 14822 480 4 wbs_dat_o[1]
port 619 nsew
rlabel metal2 s 85642 -960 85754 480 4 wbs_dat_o[20]
port 620 nsew
rlabel metal2 s 89138 -960 89250 480 4 wbs_dat_o[21]
port 621 nsew
rlabel metal2 s 92726 -960 92838 480 4 wbs_dat_o[22]
port 622 nsew
rlabel metal2 s 96222 -960 96334 480 4 wbs_dat_o[23]
port 623 nsew
rlabel metal2 s 99810 -960 99922 480 4 wbs_dat_o[24]
port 624 nsew
rlabel metal2 s 103306 -960 103418 480 4 wbs_dat_o[25]
port 625 nsew
rlabel metal2 s 106894 -960 107006 480 4 wbs_dat_o[26]
port 626 nsew
rlabel metal2 s 110482 -960 110594 480 4 wbs_dat_o[27]
port 627 nsew
rlabel metal2 s 113978 -960 114090 480 4 wbs_dat_o[28]
port 628 nsew
rlabel metal2 s 117566 -960 117678 480 4 wbs_dat_o[29]
port 629 nsew
rlabel metal2 s 19402 -960 19514 480 4 wbs_dat_o[2]
port 630 nsew
rlabel metal2 s 121062 -960 121174 480 4 wbs_dat_o[30]
port 631 nsew
rlabel metal2 s 124650 -960 124762 480 4 wbs_dat_o[31]
port 632 nsew
rlabel metal2 s 24186 -960 24298 480 4 wbs_dat_o[3]
port 633 nsew
rlabel metal2 s 28878 -960 28990 480 4 wbs_dat_o[4]
port 634 nsew
rlabel metal2 s 32374 -960 32486 480 4 wbs_dat_o[5]
port 635 nsew
rlabel metal2 s 35962 -960 36074 480 4 wbs_dat_o[6]
port 636 nsew
rlabel metal2 s 39550 -960 39662 480 4 wbs_dat_o[7]
port 637 nsew
rlabel metal2 s 43046 -960 43158 480 4 wbs_dat_o[8]
port 638 nsew
rlabel metal2 s 46634 -960 46746 480 4 wbs_dat_o[9]
port 639 nsew
rlabel metal2 s 11122 -960 11234 480 4 wbs_sel_i[0]
port 640 nsew
rlabel metal2 s 15906 -960 16018 480 4 wbs_sel_i[1]
port 641 nsew
rlabel metal2 s 20598 -960 20710 480 4 wbs_sel_i[2]
port 642 nsew
rlabel metal2 s 25290 -960 25402 480 4 wbs_sel_i[3]
port 643 nsew
rlabel metal2 s 5234 -960 5346 480 4 wbs_stb_i
port 644 nsew
rlabel metal2 s 6430 -960 6542 480 4 wbs_we_i
port 645 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
